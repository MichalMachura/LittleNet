`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
f5tp7gx95h+CqOyAvcE4MjQTXLWkp9P/nW8HtZJHi4tc1mTziWuIeDRrnBpal5FGXvsgSgyPJ8tq
Gm6v9PK22w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gGoyFZ4sUSXs5x0GDvxCxog0GJGuy51D4SpVEk1KFegmBjuFoM1TzBSvbGypYLaayppwXEafrWT7
9UbeSo8vmocgvsDFLpzIv1TtqAFgFz4Y3NgtKG+N4Rd3NUwY//zPgAix09u9r68PZqeDRnLOOimy
1/pGX18Q5otieXaX5S8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rfjUIkjlD5r14G7VxX4DWgMA8H2kEnt5KutmhJOtqzOoJMW2Mh8j0XWqosDO90KxG+H2/Fpj3J6h
QAqzA0UanjQDhWV3TsRiIiPpsVCNxfSG8AXQeN0b6+VrLHjuNVxeSdaZ2Qu2BhVza4pDeOqCz5hr
wR6lE+ZXDq9tNIvPi8Y7H0FOPlbDq3mMYoy8VHabfIEPE4U3HhUmjoNN9DZqrFSXbmVbO42yiU4q
CwoItBkkAVTcn3NSm+5LZan56i7Xa5uTiPhC83b27302oKjaKDgTgLKXolhtkhXzEgRlzIGWBWNP
1q0i0N7pCKHbA+mqsJ6TvqtkUewy+J+MnuScQQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
No8a/uY/VCLQmm9bBU8p2tnjL3IoukEo7sAkW9kgwWRbSwPnLGWYPj5947v6OJGoULPSLNR8Czlh
Mg7QGzOm+2ds8fnCTykx+vAZnnXO3FWQtNlCklimUpCkq6cQMNLv9vKc4eT+AhP6tZj+H+kLh0lY
71wafjrFSzHHGCHMBhgdGMzmCkfc+r/UuuCIwO1y4RLl+97L+mw6zxsGhwZjuyqgglpHeHKQxPbH
TdAg7SRvSbqZS40SK31KmFh1ekC7ZLTunCq/Ter82wltSFZx0BpBawnMDs8Kx+R+38Vchyu82FsH
BWtdQZb5t6D3gKd6V2mfzk/K7akkC+4/rt1YZA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cn4IgLuobbF031QXUT2JYOqXnyGu3fCw3KW3w6WZmJD+jl7RzQKGSNpPYuw55WG0UlvjJ7uQCGGb
kN3fy0Y+q3CM0x0sT7xp/H5kBUlaB764Uu/VqF1IuLUdOfkwV6JPKY8+n0En94pCEtMHLgzkhZ69
rhs7hw1jXHNjJlMNWWE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNkLq6qp1CfT5Ex2uN2F5SKzy3AS+wmUOjA1hZzgnrjIqMMUDRXqNV9nhYqYF4eeK59N00Prpe52
YyMPc7idI4WseHQmT2qpCSbclz2TxqLhIbk/fApbCBRhtBGjepAZezey3DXT7W/Ch8XQnhwADm6/
Y0HS0wn7zrfscG68qXFJdK3kGvF63zS0vf4/w0leBmklhcznxSZ33WUqupud8gcEjMFGOrUkrA8C
0w3PvOR4b8SdlHEL6u+ucPeS6eikyVVCDLegNuKRJ2co8UAf2/8MnZbjeNx99vpZIyOQv1srI9qM
i+dMbrqJ44NT0oQxMxNy0sC+L2juijjrd8Qy2w==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
exPH5U57XKLSYIN3xvaIhyakRYeMXPJjLjGBEZk5o6AmF/R1Giz5jE4r8k0b0NMJM2ZlyirJtLjX
PCu+4cKuR9gTOxVtdZI5X9LRwIbRzbfYXWeGVFHOfCPRODOCPHL8uDGuLWHtPAS2x771LdtAyyk9
m8pZYd1wLknIOtisNwvGDPiixIfuXcDzppcG7GUI40MQcFPp2pOSW1PWWtAS9S6r+6A09k9h2Aif
P2fnmr0h3W9XUzrBXQcXJ5NmxMzY31l0eioMm8cR+aKUQemlU8klYvgPX62QPPQiNgbOcQzR1Uya
c/QRMWSF65yAW4oRT7oz2/ondiPYhjyNvhkGhQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OlfxM5/8pCpX3ctYK6+3eusF5b/1nte/PXKw3/flRkYPwPbMw/RJV3S5vZF3uQbKlRqgcHND06kN
87aCljf/qnfeX2R6pfWtYCrjPwzZtPjQg3wZ+RA7bq4+rUofwUFYEn+3FGxgxI/1vbSBK9uJvfFj
IEKHKB887nRGIDrqCgUGBHmLrcYkcHjmu5ohjBXHgbJQbJXMFWAl1wj8MmFuF1cAXiyqGpuFTR+t
P1oEyQJyYTP4o5pyQwOYFQiRlYuughqi8OCU1BPZknuyAy6zE2zFDAXubmIOI1iu9ETOsaTE7nTJ
3pb/E8Z45N63XT26l0rpQ/xZOC5H071UgWBvug==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AgUK384cSbERm6osnRfkedsaBtK9MO53k/pRY9UILFf0LN/5Fu7oZqIbnXiJIGvGAdCE+5c6Bs9/
1hwEI5NyGqSNgJ433STf639rBDopG1zOTXZwxb0Q+J7UWghkNEImXmedKu4L3R4c1Tk8OwvL3jGk
HXJ1/FhxsToGiqhbzmIpmdyq3rZT8DiJMl1EVfKCE8yk2kVRV3ed9vBrdtsDjIRPzrPyx3J6bjdC
9yfewJplkOafbtoWWFcqPAlSl8fzDv8jLqSKqK8gvfvYF+BY87yvH0nbv8iqjWkff9V+AY4rF5VZ
wsnHZLzhvuOJsjLs2WxOC9ZpVgqnWxlF3twbhw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 102992)
`protect data_block
zWTyVcYIwQIb5R8CJ+T1OVHEg1ngVrkfaPGJVtX1NuFk5fYsQWKmpiIzzBCwcoHOlf0uAZrsXeY8
utAfjJWA0NjziwYEfT+wfvYvLq3REPyJtqR6V1h1SoOk6iLpKKypVlBec3Kh6lP1EK0fszCpV4ic
W1DSgI+PB+BR2gOT+meX5XyfVaSV9Hs+TOqP649hQoY1xpfNn75PIAw3cZmQaUcOuUvDtvhL5Oii
PcYyXVGxl0eXDlmiSoTUdGIh9uN1VjCE33C5uOow16TJWvCdIngeEQ2Ze3pY1FgTiWTfV3lgnGGn
U5q4dBITtCxVmXGwdeApAbepM2pyVlyqZc8KmRFk7GQRW8usW5gfl7xEOyakDJpUTYGTy92Zl/8I
ifzftHRNmXHU5g7/1QY3Gg0zdagtKxQywiVNa4kEfJM4nYCkXwO23yeBt4MymdmROloiq9ELG1zz
zocEbHm62JdcNGjYRglEzUVqt6nEXHPEWQgVAiN8gWSfrzkQNHxeWmdv3rlSU0dWouhtt6+oQihT
0wHP0SJfZOZRjZY/VBc5XnxoTV7yQfWD5xzZOzxHTHZ6kItowccmyzHvPndze9XxUddIH8Ybmwyz
LS11br62yOKX35TQMS/EWG3jS3dFQjZmwr8kT50zGcVVPDT/os5EVPQxvnvXekkCvODaoG+eOtIi
S3TbkK2EpOc9LGphp0OY5sInn+lniq/ElfqRdMjiktdSVGyvxj0HcGDhoIFe3PbMHW9dnmnE98yh
PczrguMfdysqBHeaSdllzT8d0u4AkcZnYJx6BWK6RvyLwm/9gistidl/1lQQQsAzmeLtFO4MvJvB
ibFnNxYQCI5/RTBzTjADv7yhjzFVpo631RJGXUopyajXkrT8dFyxC2+AzzWOw4n3Rgh/+GOqqigz
LYv9HfSvf9GwJ7zNastOjFqDRScPPEeHgEV4a3jVgqUxyMGczfT2kgOGebZaxCpMhd+NZbR0wjfD
vkJdKKBdpn5PDJsXhhN6wqPLslhL1BfA420jFTRd8w98kThbXpO8cyf/YA50H7x12VJedYv/nepU
rohncy2BBrkB01sqXGce3T8P5yOyWlrdbMLQIUqLfWqCFpJLrmDCf2+MOIKgKuwWT/f3q6R7ztbQ
zcMGpDJq0D66n6oRNMhnnkDtkHecf5i8O16Lm2KDYrgqC45m2/S8qIw4mnZm8oa8V3BOuzvxYupp
gmaGNk6+nG54bHulmQy+vNN5RHB4nn1vkdVrQlnB678ROz+fKaAZofdncuYYo5heIzSK1/nEP+yu
HEuvdmq9D7/kt/piWnqFURjTi69Tx34K7U35UUyUpri+n9l3SeXnubuPPxNAck23lLqHcKM7S4EK
gVy7c5vyhy0+lBRhN4HrQOx+yN1i7fxohzJlKyKUSEBbhHxYb2VrWpfAatuGfGLajkpvNuDbO2mJ
IZhEcbFpIzYj6h4QoKRrzbtnJoh0CThAnS6koqj+5a2iOi5xSZSXtcg5GjgXqQVhVR3yYBhMLohB
rDQWmFgf3Y7qB/GIgrMnoW0ICNKrjCgx8Y7MPujhj1OEfwcEMsVicvYO/+2WbSbdRhJrg2GBXlv9
yz95H9dnbF5bgxcwXsWdOoAK8Q5stxttcug4nGruJJ6H5jdtaQoRrf++1wXNsrk6LVmHeFO1FN/8
80TrHmL4r1fW/BujLHieDSZrrMsb6EG7K8GkYmVQXRuKTdABeFcvdIzQ7xnNduDhAWWNXgF3zdQL
ZNu5aa+caHyZJA9BmR83JtKep93m+Hqo7pxu4d3wOOkmRDFQFfSmE4FcEDnKUrXHWF8ukRA1Cj8v
l4UnGIQVBC7npA0CcxdOa2X1TaiK8r1p4JfiKCJUDR1aZvqyzeGErlctkSzljo33lVVV0TKUdiH1
GZOfg/MfdneDP0GwFn0SWUukvy/s5++mrm2VLhGk6/a/tsdhzCY8BN1TJ53jUVyzmFaAo3NG+wxH
mBstVysKLVW7c88Q4iL8RjYgIPxWz5zhckzr+E+qsIok5YNmcNXHmdsY3drYq5AcKGfw2kFTWfKO
hdyg3fAbQ3QpSRwvJrbb82gMszJUgppW2/lEqqhuvfrTS7kNbCqmdI4WVbwlvKu9LV4D1kixrvRN
YgtCHmCTHmiPX99gKQzXm+Y/31oqaB0eIE7TUA98QDnyK3oo9UkXAr4R1CuvFmATTSg0HuBk3CgX
zFBzj9zgfa9ara6w24LdCR0TIayEfJOPy2BCRyvpKId+WlBcmTWz6JbJD0P11nugedat+MEcSrG6
uQ2amWM7QtGiHnlhviJX06nPWknmpPzlo+HSG6yQHQPDWFbZv17kxkgdD8IiUJ3QURDjLSRvW5ER
aD6bmP7UopXy1/KZLzsKUfZIeUjuOFD0i+U2udNIDBYA2eZBTQcQ7Eu6RiHcCwptQqLxlC+8cBDX
usRLpOF4ArdVtV47QnS3+dYY8HrmylED8JAe9el8N0i2yaHdszIIo8XKZjsIeGHmQMOgFpz/ohjq
tfWvXwMOU2eCBvgK+io5XIKJ80+ujt3kokAyRujlyWNIDRKsib1AYdCCGHSuQ/2xHnjx8LxktGPb
6sX8XKAgVewUBX+GF4AGzXfewRW23EfgpJ4OWPa8803UrcS12LoQkx2tqffivygXGRRRKRWN79Fy
TmI6vHgws6RJaEG1G4EOtjQw6nOtCaYASDdmKbnIgQxv7lkJIkkrqwOpEnAnmcVSw4QbhHp6cq93
yVg9mCu2FtRP49AS2NYC60c4Kqlf909Gr54Ord783hs5PJT+A3mSQIMgNPsnYzMcPpPZdIyF+Uee
iVXPrbeiAee3L+vdyrzfuTSqFRe7XQXhWprdLqIL9dIt3242JWYJYmof6NWTDq9UWPQffxmgxFr5
NiOD1mAoJN40QqwiqS0u6rdkYcRgGQLFsKxAZUw+st1kkcgrDNYMG17SO5/5Vog5ZyzF96Lm6bDJ
0k65nz2CR5SeeUUFj4Q7G9fAw4RrGC8lgDklJqPAE/PwDQHm3D1PO+vl9ig+5K4Pp7DPSO+O+nlA
mbnUTREZSHnUu6nKjZrdnqQ/hyHTfYVdbCltxEcx9CnuZBP9HdVbQG8XtBygClDthidOOi5g0Tbz
SO2aU5apP1vJUl45D6kxdD27ojB+hWXw3lelb5AmAEbJ48t2A8PDaGtMX28ap7+HyL69TyB7sEZk
0LuWqmjSfb4bBFtZw7GVqNydKECpkFammvQDZS7NOlqeVspgBPmeMGO0oznojFtgztn/fhmWDIFq
3A2uxf6z/yK6D3Shd+78+M1QleUJ4Hho3F+fhU/DZGpMgsUvVk7wzTb45JTX0tCF4DVZ7RLzgn8N
CPnV64tYDaLEO23vgMlE+eicK1MryziYDSHYCTrnLEADOZDR6p1bM8JEUI1iXknqa5zW7s2BQyWj
UKUSzikm7+zB3IRKR9cSpkQSMUcORQHH0sywC31yZhv9eA6AknKhDBWUUgrQoM6LVUErNWh22sit
2ZJXPcFUf0Qt5tNR8uJDUa7o3UNC/HDBGqCamwSjQOLTT6DwszF5ae7Q6MfLkObLAxBEj6hHb0lB
RILuCbO2XZIuomspSPYAAW950XCkg0fYcG+8m8Uy3IOc7bv/OTEYmIDTPMWqqclipLMHBXeMcz/a
2MrfIV0mMsKrc3FA9jMEztLHjjuoAziO+nwCoQZSKTmRmK449iWRXOOr7bjcmazqa73ZLvsnF35U
suhUu67kNbl0Btpr8NITv6k/XG6jlx0PF9bt6gPFgIBqROO5mliIQ/1Tc89LLi7/Zu699S0vxkrz
7FKpKHunCjDQYIk/IHgwF2H43JG5GTQsjnBHVxK5cQuIVWtoAbvAEndj0zMLzpx59/2Bg+jvDWRy
UenWyODV+wkRSEdYrSQuExlZWdsqU6ZmqN/WtnYxpfNVJUlXdoW3sR4ijiWU2rpcw4UgrK/olgqN
g/vOKCwUD92mWaJooxzzXo0ItdEXWBAe1GAl7mc7NueHVeI3fIgAruLYWec+KnK1D3pWVCKnV5nR
x18FOpqOjU27/4cTqnks/sQ9Ojtaz+T2IO/5Ei/obiFGaprT8prD8LQHAc1q1mQbZfGmminFYAU/
pWsZ+hNnqW3mHB79JNR8N9aQ1Ej+4xhlaNf+DDAV+ynLuMS6Qv8fnsvLVN9huChxpok4hml2KyHw
Ux7PjFHlzcxn/qZGBSoEyrl2y/yFEZdjPh/ASXKCTN+VIQZEiwZV/MM0FDvPsiCnFL2u7QzUORy7
rCFq1Aisb8NgWHSZzGyjnmSqXim2NVNepMHeAOGyxr/E8MZQof6npk3xKCyxt90+qZAj5D3FzohG
ibu+ZktEbRnYFVqF1HWsMFswOq3vgjTOopCcyCszShwErAJSgVTBHs/QzdMk3n4xO4+0y5NZvWFi
8dHTpwf5tIifiU7WtxpFsqe44yzWC3crpSxlkLJQcZlwpyHxckEgbEKJc9AbJ6YGu6e/e5xe38OR
Ejv6ZPJm2iSYjxeVJ1bYhR6h+m60lbX9M4iZBCf1G7kUXGTmSvo3HnrajCPVv6tmqqLuhaQn6k/c
eoWjMrEdvWAdq06awCVuX/cpMk7LjS5+4rrqHhyqfBlnhNSWqErPO6TD4jy7vsjWnnC3A8Ki8urs
7Cl5y+5GMdQ8Cr6bqjs5eMd0Ja0FlxEglQY2SPI1Qc7+3K6/eMofokr/ZY3b5a0E/L9rfXzHejeQ
PHLE7AkO5Z7PZd9bNVpljf/MjpDdU8jhmxgjwNp5emfw/RzXjgoDztKuyr9LRAS5Je8Skhm68pR9
iFZCv2kfFUJGCCfOfEFxItLgYH9SCmukD8ABFOi2MRBchWHbgwKfG8zj+m7Hyccg6SRzqOrkf7ap
vfpO2UZZMEefQXpke+pDeYppj3dtxcwhQVK4ENix8MXyAadYL3kK/fkEC5IeLAgLe3gNgawmsS5K
rOqmWAGUvXjJ8AYyfcRuDlqBaqxSu7D00UC2v65akJdGlBspX4wUDBqhjTHZCHng6/DFzaUtUdWS
NPfBuVqzK5YVTqrtxbYiBsbBaRCOdCfXpGg6ipjXmu2/V/iwAsX2WHT40Dp5z3g/cd5ndwj1RKEs
W7DOVNl5QmCUWa5TKJaEo5DV3+HpjG2ucGv6N+sczSGAb8AmrrvamYFSDWXgsnRy1S+Yqmx4u56A
BKDPJkr42cDgjGIT34Kt5TDiDPAhgS7WZDdNbz/bQFDyj2BUXmcvkuHk2RHmYSaxtsS2kA10D1is
f/G6L5mwD4P28inVE9bAbDXeuyg1sJ4UGWNO7MJd1ow1fPnpV+ZrBWqKxuRj+nONFuuwgEaNe57y
NzrLCUi1ZJNN49tBBWC5Amjkm+d9QW6qmIskil/sfh8rLXw5ilVDqzckQJun2LUjavfGlrz89szZ
pNTckb/ZNiTS9plLKSO2O+IUMcQn/z5JiUrDguV0weCoW84OZohgLZLKATDQxuHctFsnuubk46WN
j0RHuKBPclIassTgvehaKa9DrrwwAnU14H1Cu4xbdS7Z0Hsc9ErM+LXPfXb8g4OZMUNorsAznCns
VAHvnJSDQZYCXTu8IPmtdAGmTN5mLN68F1ZhYSCuME/sVHOtwBV7xWc1yW9GWhzaRnyiWlsN71SK
A1bE1ui1qls7IpSYSvRUdarTQzMr8MkNuXjHL8OJ4X7o8f9pQL4bWMYt7kTjk/bVrz/okb14djyC
/9spgHPTzbwwKaTlOC96K7HiTcObmifQ70IQh0DFm8Jg3jg6e1+Axe0m/LxIKOHf7itW2ypfofGQ
xDNtS9GE1RxPKleIhlCzABqk/otvidCwMbo5r4fP1ajlq4UjX2kRFM3sJSzrpTKcrm7GUIQs/8b8
TNDxa/8+WqxC+pl5JgykXvgXZ5faTXYoJp6/nPpVZYUY4A/D0rIT8xyoJ3+S2Dx9zNdTZtg0vu4/
DVSEM1+csW1qOSAX/a+QawCdN9eUPU8zPM/bgXYfEC44p+6pwlXPeseUb1O5e82m5tnZGLwLl2Pl
vl+Lr/1NEtTYuDiW7/oR7cnCg7lPad/5uA2kzMRJj19StfCSo3Zi4CrfUPl6OGZKct80oDlOSDqX
Nl3opd4F2zQcCpklHCUFrxtTdHqNljvMnYaMLfVB93QVsfV7hd9gMZr87FemFuar9PzGKsHbvHmq
4DaeWPCuSnAFiJ4MWsYkgeS4PJbpGLkxHOfm4PxEY5z3hslHkGBoyB0hZBa/saSXGnpgmVyOioEJ
099WfVdlLzC0n81O0SFomy4kis4T8PcBazCxWWwocjEJKWDo1T3INHYkPt90/gyvfnoSo0nG7dOk
nxu4LBM2ruc9Ezs1hOazl+GX7TLfA5kTBk2GgzPYF3KzMpwDV+6ZQtKff9xFKNGmyVAYbPMw3Xtf
jOEtihkyF8KihuWZFM9aVFeyE/N9GWizstxoroYEg1zKSP2nUrOOw6S1zD7BF9yCt7Bmvnu+PHwE
1++P1il925O1XyszPHtbQeDn8qadtsWxB62ULPMcWG/elnwcQjTIztjWM5b8oSBBPmEIfgSd4nJ0
Hm2rK3UtBm91asnI63JfWX3A3/xUy+GamJmFv7Q5QbBdN8DbC0WRQ1c7eonPU6lDoHgEJVZuL7eq
GofHfdnOVsMv0ZvForx+QDVjRsb8A9ttfqKYiOL0GVAeewkT6st/ItKbQKOHZPG4DQhaWYQoIQ94
mNt8cpcVG6ceeO+Tvx7uZNNL/EURCgiOu4bnJHQdyToVdP87IBK1J2UOdNElJmzAlQwK71fw6P30
eQJpCZ3BeTVsjsLxGSaZC+lTZ/evF82IERa8+NlDhppI4hmRfldmBo/YMhB9iisPzH8xG2WpmIcR
oPzlaTSWjYD3e/NhWKl0CKHr2F9Y84SiFCKMlaz7eMiU6MtbnnhUjtDOTxPu+jiq+VoGIGiQT3eA
TZmBZPwgCr6hmE/JDrO9317DgnXVYHoG8ZItDxWLVQ3AM+hR2vn5ShyMzGioZFwQ0knY+uWiS+66
iZOwDFTdvdKPU9yNvW9mkbW+0//CrO6o5/GEDDK8J17oBFyWhgZZRuxQeXU3Xl6wlDwjjq57MnkF
uwcyrrUlj7EsJSS2IhcPb4v2MR7FN81T8VtOPeu87NqdRhnD95kmbmH8mqmPBwMTQCb9r7uDfx5o
qXGPbRStaJiyAkudlKvYz53Udk7bOPevXHb0p13//n4jNcwNyFdI6aemmQBV4Ia0cMXNNHl7SNnl
DnV100NF+woZ34RrAgZnrFJW+zWEhrwEWujcmCDD5o2iu43USH2ZjLVv0TSgih61mutTkuo3G8qx
A8JuzyeU0NDKB2Qqm7oFFio9WZcXhKxbMooNAKS8+kquAcIdHvqSSCoIazw1y003a3mNCCB+Teqh
QxaY7dGBV5+wIgIGDChzeDRVeUZlCE1vEKAgJOUwYM37QhNPjmvl57cDXkKBOo0S5AKbSCO1ZSE6
0R9WFh9UIy90lrqv3gy14LrVFJcSHvjj13hrwYgQokVzH+ibg3z68MfFsXjQwdV3QNF4QB1QOlD7
YMMNQR6a2PNw74k7vX+n+ayY6B33s3YPn+BzMRMzKOx1GukorjVqS9mUmBLRFwJU4g1UbbNJbQg3
hy6UHmI1Kq2GKu8ySVrme3FWFMNvpIkr1yzZCBZuP28J9FYINNfwXgoEGJ35DzWS6F0PnJiJzt05
s1jmhmGsBFYU/YRxKe9insRD5LOS4o9byMQ+ivLd6iKW2KwdwgWuFIcN9iy6q1h9YwpjvUQH0Iw6
nNXzIEtA5IEyePIwu1FBrRlKYV3Hwey+rzLKvmoHbDgcrUZOyN7OGEKuaixVSJ6yulsVD7nM8wMP
1ZGu4XBrYsYbTCzlU6L+Okmk1jtdTnpBYnj3nDCyRBI4kTndadC98+3e9/15iohFuKfA8hmz/NTJ
Bo1ZRgkdpR6NRNLCMu9fGgpYfIYEF9BS0fxfikdea3FF1zdNBLtaGLmV6aNONXXl44vhlOZelsL1
gqiHi5UGKX67a4hQWCQvvPMLgTjNJEeqWUZCKoOsdsNnJddwbxreFW6gHE3hCl2kLXFv/A7D3mmK
cQmmIgaqdQf49ykksr4YCggVOjcoyUHNpA5TJv9B0NGhqT10KIMUnef4ToLXZrNMGNSunxC1YJ9c
DqPUkMm9kRgKNAVt8HDaUfd+YEG2QskEQF1ueBobnKXcvk8R6fSftGcItYbf27q2cjK4kmlKmqAe
JeF71DGjwjEBqhIFfG0MWWFoSxaEBl+fdC01IXVJ8Lz+BeeCYDAmVzLbFShwO0VS3J6s6pso6lv+
qAK/sT8fmOU39urA8R9vTUt6f6CLGSi6PQTy7ef3oMbmjn4NYcfQdBMeYEFrtZvH0wqZf7pPa3bY
DddEsfEYzuJjPDoQSuGmdDo3WlIG+vPgQfnEOEM9COq37dXARffbjzHVaXYeTvEdVNPZWGRd6xuu
gKCWLw3ZKu9jqH86rAxX1n0jRm0Hq9PWut0cwBom7DenfUIljbXnSjj3kEVm4z5G2OFozXv88Ku2
J0CHgjt9lhuxyN8Wv0PO2+l+RCB4E2yemlSdYPOo2Sw6I8+psXq+fYGkTDbpllS+PZv87rw10fRs
awb7USopHPeq85PaAbq8AtYNVAe5oAdkaV7LQhunfejYlviaZr+IJMH8goU7eaC+yPoB9DopzQHs
/aZ7oHzmfiT+5nFoc/+udS+gT6TdSwA2HKGtHq4JZiqbB0CSEKnznbYNPF7jHEQXD3PO9rltJojm
fM0Cswz25zjOK6ov79nruRBgCtFh0JEDEGpWwCTe+Ldos2qTeMCLWwT0QJ0ep5e9cuSAOVjMAS03
8PgRNQu6lroSMR4kmuAum22lamDD4wNHrHgCixB98M6NQmVVcn4DSSg3OUVxHTUqU+z6sXKDy3V0
3HtqEiQ3/Z8A6u9um0RZ6b5BRh13QbGn1Dn7OLd5uo/TGkve7fAkXs9ACvigO/2aPXoJGt7j+KV8
kgq1lvaz93rEbWu5HDG04rKwr7KAwHmGmRdG2ELu6CgiTVOAKXIO0grqhb9iIk/zGe6T0Kzz9mMM
2uahE+SPN1L5qlYKwvtGn32QsjuY+75yCrcnMil+zpFlvmp8v2l5s3yyIxiWxo9H5ckOpSFYWncQ
OHvQBrD5wTQAFTMoTvXq/4FdPMELseNcYuJFp72yqh1Wdv18MLpCf5IXgCiQiBopWCynNnAKNqxX
HAaKIMZBRxf5ejmb4+vEbjAVNtJXLVfseoy9U92L4Fj4tIs7Z4uSsC5yH0d3vH4To4rY1gWu5SUM
h28NfsirUHK/Y3P1xfT/xscYL9zKcqmhaaSQN/HrGdXl//ebxV6hmH8dGu+hnLo5C5gWpllWOwXj
BfcpTxSOrORMBn5CUXMu3KROoZSatm0r2NxR5VTfo2PzWfNd4CzFPuSxvy+dNMi4ewwXvhHwMlI6
+zAl30Is1pjrdAwQJnj9asC8PPEzdZ0gSCiddTRRxOT3wPmz4CnlhbKdWbCOoU9RsObhhsw2y47z
u6MthasQuexE7wJqS2Abey7+ynHhyIkze3Ye1RDOFwhy1gYH6yxOa7mNeT+pvQfwiLCMYnMBgncg
M7FcVr2BrFwsn6qBZWI5DPpneL9pGi+kv1RKNiroUjAbv7/xgoXYKsVZeg5J/jztZCPndr620fxb
obBHNOU1b+mNeMAmwjmSR+hPdHxvHO1pksl5ev/jC3wFdEnXlwf6Eo730rCft/5l2VfjW98m2//a
2HasajE2cq/Ig1WN4rdwl5/7fQQQrreSa8JQA1h5HamJ5IVs1aIz4NM2DIvZHbOdI4HUD3CodmQh
eAVCS3H9NfUAid+FTVytk8UBRYhlRt0Z/bFTZcP4tlrqKazhRit2yrk6T6NoV3WoV2H49fu5VnwL
SldNWslAm4oh84i2unt5xwLC3PJuqLfm5cZjds42d61drh6wCPUn894HpvJgkpWruc3rW835xSBi
HKg7VOM+m9OqlODNywsn5kiyQin4AVkZm1ngtdjZRXCwDmDrnyqYOoKJHFTKjSE51n66ZhstO7iN
P0/+YXJPodvLOkN7YRLCvTwE1ZBTH+JjuwiuIvtuATQfPLyXatSbfbAq5kvXU3USQZJqp8H9vkda
f1aUlenqXmutSbRHpVOa/+m2gSEO07f9azxPRh4ZU9OBK0pqCRzoEaQhqBzfu1W+8MtFvOIcsw1g
/UyY64b5U5IBcHpSO/cd7d8hy3c2MQ6jIxcuJEzaUh/zMrrkSjAo0ButZqWIagesdCmbCx//aYpz
dKzyGp5jV1iJLK+713Ih9DJsYC7FebgQpPfHFNQT00CMZWrltPvf+TNIJozYx16Xhf7T/cw1Ngzn
AThE9cNTKgrxs5Ac8yWqGImYZdz6NCur/VSJIhlS0XFE+5Lc/x7d4QNht6joO2KMcsd5dyNkyvxQ
Cu2v6fd9l0DvwzoNWCd8h3WxQbqAC4J9XZ+KZalKUwsRMANcQmgO63vhuriKEEQ3o8EnDf60pNe6
4rPK0mEi7V2JekG51S82btIwhFUdpgmwqJNbPzXMWND3iA+zwZ5qSFMF2gjlisSefdCUG6g57wSV
0ZIB0poIOhVX5/t9DQhwfD8nIKhPrjH6Q3EWbTZ4fdfXPhG8xW3EKx5RdUGqQe1r3cShuJUFuJHk
D8+c/raDCEhYuitjuAwezLPaHeB+VDyI8YLXpgirU64zQR+NmD1cfQmkmX5uTSqefcgyji6CLKgO
lel9nGgu1trHYw68xeeq8WZc1V6Xa17ppUkW8+SegsxBkt1RLizzRsE+4VEOGVh5MpjBIAF7kbiI
U7VLePGob4yBUTBrKkuNu9o7QpIki5RxfuIFXPmbf+bHk6YuqdCpi3agyXOJYCcDE9Fm6ymbRlte
Zxhy1tzCfeCSma3HnWHjNoLukX3SFCmw7Bgf6hQNB0rSlVB4/+EJL4+KSNFNH5P2XUMk5B/RAhuX
3LxJj30srV9C3onmtaaHjJiA94zpC0V3uCTDmceKURNk9ehJRE5m5xJRrcmCt/pB+S8IqV3UXTt5
4HpATpw7yf06xKDkU6i6d1rotgNp3ckHqEgqTafsW3B9sP7C3hBuCP3peIpUzuKF/wkBHrzdj2CE
PMIvB6jZhtCbqJM3x1dZ+F3GMSTFU8mg6VUCNx/567jEpXr6v3INKBImHS9qG5GtmTXs6xHeiQEO
8LB/I5Sr7SzyOjI1RpHdWhFu3Z/g8+6oQUNf61lE9jVL5p6DC0x/0v8jC9NKy5Vy8wXcFHFDYtek
kFmAniiZuQgOZtaMulVEYBF7Tq7sEN9JEEG3nIrCzmVuvIBAgIa6uAcH1GYefC3kWBO1bhjOHhQj
fypg2SJz//fS5vStof+A+FwUqkTRsO9FUJrxWiWbR9E1D7bVgBw+dTbTo4q8sMRNhVZovx+ahCTu
9vYA6YD9qol9mWda9e/t9XCKDXgOefjejcJ4bABhjfqulTj3m223Azj5dzkMDz9srCU2rykQBGPt
WDBVb02HPLYygTnPR1l6uvQ6HkUuNsQcRfTNekLVGFaks5l1Jjq8jO5lBBgEwjxDfHwWfgJeOOxh
+y7GiQjYS++YKdJ5Bi1Sq7JhduLnlIyx7fWS0LYqri4CLDizHSJBXdNmUrSn1i2NbBl9SSVwsbuo
mhwGKrTQNxnoJVEIGQj2ftGhBf6g5XEqvfY9j0/w+12HCgcqjW+RDnqEUm1HgqKQ25JbaZtwtZ79
f91RZD0xCPzi0fWW5lV/rQPf6rv/UMyH4/5pdUd3NhTLoYMVre5yZzbJQFFNrv1DZZwZ/3HFPN9x
jYHNYl+f6MsG/5Cn8qlLKK6Tcl6CXxPVyZux8vMm0iZ4rRzZgp0UZvSoyslBvhqkwM8YPYjLjTTg
8TCHMw6vNkkPBSsKrI087BiYRoWz2WOxW+6N2T7Yobns3AKplCbm6+lcNv6kIvF+B/TCurUieNqe
bQnrQ0Dib7YKjVXxXtoNifEDwyVQnMpIIWI1ldG1IrX0WA7r9RSjigl66S1A90Vt9BEJFquey1fh
WP8eg9bBBd2cFZcpkoC7ApeEQh8b4kb63O/8ImDk3H2t5OxsqRTtLmg6uY4VIfKe2PDy2N0R2TnQ
+M41FSzr/Z2IgsDK26a9ms57lCdoiDyWlwQiQVmreG8ZlRh8LjjvTiOcNZAoU8NE13GnAMBPSgqX
rXYGwpmFXlYyLK6MewRN/eJBMuZ/jI/RhrueJ64kyN9ucfAdBAdaNfI/8P9d6c1DVBcx4fjXKO4B
d0/dRCYeK/vwsSwq4zgZelxjxHa8DDOT4k5KipmHmjkA8VLKKUyXwHzGXHFr+zL4hl5DnRVIPkvf
WMB9IfRJqqEUcEYv3MLl1pCXTJOZpkX6VCiTh/2y3iA6EiEkleoSmr+asV58H0YRCaKUosOF2B2b
DNgsrEjHVIYro8rQk8QNjZXqi6l0fzJ1yTU5E8Brw5wZscKMaX/QN/uzX1Rh54obtHTJcybuUYLC
knfL0L7rroZo/cEVTwEP91mSyzXgD26OhphcNLpj2zvpsON42mFNvyljhIuR5bEyBDbJFyS7cTRQ
Krzk7rCEHno6H1ltz4jDx8peHkEC3vc3FnX/GHmaoKAFeFaGABi051QQy8J6QXMs3FqWlFdhGSvP
GFvnkBzAz4Jvm1BxjQ76OrrQsuFzjf71D1yCcYmSlQbFDjgbtEg7r04y8mNZK++26jeyEswTT9DZ
BzbTuGU08jvby+5KbQ/om2dE0CMuriQzoazHJ4ZVW64I9M5MGQvXUVdM80t7h0m5f/8RRH5LdPO/
D7CiHE18tuTALHqsCHO4mQ3UPbu/d5QkWtCezGS4MYWarKJavB27eCqs/6LUZo1SMUJobRQ/mb5o
pFQ9Khs0mf/RYONf4aG+wrUueTQwllimdS35I0B5SDHmbBajdO/xWbKZkzC2DOsbSniWP1To+Ab0
2vO7BrTcFSIF5g8HfHDVa3OqhQnZCSf5CWjH5Zj3qwMQWOXwDirz3VWxWnPOx9fpdZtIpEYiFsVJ
xcBlhE1Dr8ymyGg5c80+9L7DyNzbiiANdJa0fu3u+LYZZW6ugVoo+ztE/YhaP1UNiZIWEm3Pcq+E
B3LVOZ4S7PcEmY8uGtwmN2g/wV1EjMYdo+2dG+1fERMGvTnIHlb/5uNTE3odVqqqJoNvAcvmeAGN
wHD3MjLPqjegf/zg6HCTqqensk30VpHo2JU0ZhDO0NMjIZOJPUoQPG2/NdPpTXTsdHQphyEd1H1y
/g0PJ7TAlFRXZUoz7RMCBJ8H0kQa1c/1z7OcEvKps6k+KLhKubDT21lHAAirnp1MXjJHJLbjCN5U
OaE1zV2i+cDvDBuCAjAh8bnamPRZpq1pl+phfYSfKlSBfXaXhdI/Ohb+LLsCycBrYEini1NmgJ9F
3JlUb54yym39tDCOb13wPjzrg6pdF2GMrNXNC3Xj4c66xTqq/i6k4tXA83phocXN9Rx8xjmZCC66
1Ljt15VlAgFGe8QqkE/A5+/r29ze/0GBGvHiufyBRmgJou4ZbIwRzniQeAzSMHuAB0YDVleg0U/m
mr0FA67BnoKIRuharXFCH4fOaHqX+MAk/4IIkTDv51L8gj6sn+0rI6oiKxWkFserAnspfnH2UWHp
Yo+Vgbx9XmzUJzJ7Gv1EtMsxiC5ynS6aLT7OqYjwKhqjZInBxJ3G23uGNGXdGQCAV2AWKck6kwUH
SUF2w1k+DsGlK2HyewiM6h0bi3ScHq2rYRKR8lu6hezBPxJzDmb4EGb65QDCqx9GWD3AY+mRO7Gl
/Y6EF5WgfThFbDUcQecFPSl1/52iSmScb9IielDfCNUZbl1Uo82tM6QyIhI7QH9Pk3fnuIp1S9ko
qlDwSY4xm4Y6p9cTf902Jw0pDVyMfRp3WWRIqpHVlPDFo5hWyQ//4QkAtlmJFFodDlnKZsXlltCh
Bp6hXA0S/8RH8jGq+hHV5ku6vINjHVpYVzFBV85qHvKKA2W7uzpc74gM2RgVnCsuTLqYtJOk+Rc7
BMJ9KX7vmej/RrzKrDct468r9Nq0MsNXI/dvw4HI69FzenFz8cPgin/UxvMv64DCuBkw9QGPUsxf
qhCZxW2E5Qq22v2NTCagZ3VXwHp4wZglU/XgHwBq+WOhPW8vAb9YCbjc3nCoDftNMw/2xdonDADi
XFiH3Mlv8bM4+tfo0FxJiLiY+iSD4NaRXN6pcToC06B0NrGWw7g/0wnGkD8q2vUnixbl3YMIwXYK
eKrjXGyMmoK46J/oAhy9JrAnl8++uGA76WCnf5XxrP+H/BXvoF6pd7yEj46aXzQXxgnkCPNZDOHd
HMSGRMbjlLbZZnJlD3jMGoiCOOZLmq/qXrwOYIvQMWopOprPRtJ0EPxx7lTtANp/bjd+rrYqJdzW
ocTESuHHlgM/HRa1Jb/B2hLljbSajUpwDq7ouDju0gdsRxyI4YBPneyglc7YtyL50WYsiq51zlBu
NQr9WeEmJuFK2e2IDkiiM6SyeTSO9npmeTPznR3vLmf/a3ZxznqAKKlolSWuznnLOao39VMm2XXv
Axzwb6JHtkXgebx9JEIUVXJ0FGU79NjVmuzNw4Dtv6+aV8SUT36DTVnyrwaxOuXoZQnVCP/NLy4O
9igaqB0N1CYBcxfAPESMFSdzmhLiaVN6XWmxbHFsvTMgdbvs6fguLP9VeCyidkA471usYoxWd+4T
o1qMaCiaVtAvMGKdWfqi0ufwfBW63apLxDaAlc43CVcUQMEB3cuRMRrXyoqeqSWvONkaCCPEKl9r
MByRL1rTt21RtEvzUIt6ocaSUkCNkueJ2NoCqtiQkyV6a2qY4Plp5hmdCSA7PBMyZL9O8GfbwOFl
6424rhlxFj7S+1FkozDs0hvDkl4AnbgctRupv5V9ORF/IWCXz10US4tOeoi5rg91gC2VaveTyGbV
rzEgG8bkH6G9LBki6rZ8BNq12QyPXwfZ1OEivH/atesihh+9DEkBHBFnqf2SzjypL6GOXLkQJTLx
hqjS9fUxGt4M0/dKa0JlLjYACFdbTMUMrJPFr4dUEwKrrocUAcNn4rn81RnKB7JMYLQWa7O5Txtu
iJdvzbeDfa//z66onCuxYbVKbb+DEOt+lyciePZIwhrdE/0i2/qLDmGTqMAEkMeVLbFYQAT/9i/E
mZJhoPAsJ2kvc6/q7p/Q7Scfs2+JmY2npd8DsnP0kXGNJ0xfxxinht1lWtIHkNbPIZyvr+kapXuq
EgabgiPpG/AqyY44vt0OYFcj7U1+hjN71fx86mNLs2EaQiKOJ9CYQ0VrBA9wLnAlremVDSor0KX0
NvTtsdEgzFcJ31ZYLx7mZA4zVJp0awjrdykzffNNxoldcxVPCBnm5d7xUbMx6kQiHAV8yga3YOZx
r+WIot7zfHC1nVsLUowJ0bMHM2nm3z8aFvxwLsYQi23woqd9C2dfowFMxemFrToZfBgxJHR42nJ1
oJ2VTjf1DlobiprqgMwUh1Vh6MzkvqJZEInPdQ+/xAbeYI2LVJobWEaM/B3wn9KMVKRAgEAfJSE0
huG0Ru4+VuByiM2On2U6EbtahDRD0x2+X4RxFhSZFbzijaBZOtPRgWhTOSwJxDU5dCvYIL7L5tjf
DNHwXBFu0WCwBLU0r59Pzu39L2flSdysVQk94NISip1NyhP5lQHNrXx8zRpBKZA2NjqMffMhmAUH
Jl7OzU3xk/pWR0MQ0yhQ58uRZWvP74cnFXQ+aMQ/df/5OSG4jCr5Ha/2J0+teIY7VTLy+vsFgvsB
nUC904c0ehdvcM8qBtA+5YXAPMzd/JJZbZrcEzrJJpshiptSsjyO/96MLz4mADbRVHM3VZieBSrc
rRvbwcL232kY/MCKBkTdnYrvmNU86a0a9JIaODKVqFsSKxgWFatzLLmS//JfALUw7OqSyGqInTRH
3Sp6NLW/0yzvs3q7t089rp4frukxnHBpyqfFNcJbP4SmBYZRV0gUHWV4w/gVXKlb2GtY26K7Ekbc
KMNlTjNS9iZ/jYUOBJM3FGd3XzPP7qBFaS+SqNj6CLJpCoxk3IghyjR7H59F2kzflf5iu/1GJDs5
1apkuAbdEzPK0rzRbVIrpOL0LA73u+CcbExBtvR066Qhq6cmzl2LH3Q0ARizdkcALVc0mxkMR1ke
6a58MTKZSUO4JGclbcyMil6CRJoYFlQUcxqmO+Y15/w8Iez63ESsLPMGfri0vbfwgQgla6HJuYCo
lhmT37thiJO+yGkK/dCDmrRJ+Z7d8sUmoP2TcjcLU/y5seOuDXu72az8Df+HO7vobs0asWCtscCB
PtXwelaYIB6s8POVGrhwmqO/ucPBAtdT3zDcbgJmGczu+6rlt6tcfijUeTrgPe6nXW6tTyMybOCY
YNRzD94SwrkkkhE5iVCJ8/Y4192U5rEIJ9B1dNano+SPCCMchsDHK+owkKp+GowdAs8OI3ZQZttW
prsmkjqSC6KsIjLOSDmtYD43HVSbKnsHKjg83qKTECv9s+dZOjgQ0bvhJHIMb8QBjtRztvqKVM8e
9PFE61Mal/6sOR0cnyYQ35HM2ef5cKdcfPoDEyuLdips0BxQXc0A6QR2Yl8tTopX+wwqkRqvoHgH
BCUT7hUuP9HVuMxuFKs69fGasnunVPlPMaKucsZHmy65phSWgn+F+eRc/91/29KI/FGEzb+Oe87c
0mcup+4mIeA/ffZJZuZ4V4EAMjHxjsXb8tgPnPwRkIqKfDdZ6ms/RmSR2YPpiAF8o0nQ5oyoJ1nt
zAI5EFophQB/kx5WcUSy3IJXUm4M6TbuWGN9WnZKYT1H5EQWzkIqvbcDeWxm+8qmzkPtp6Bi6r1/
gKnKEtobrhw2ryQM+PguholKcPdhaDw3jl/DMQ3R/zzK9aOjlDwZPBDP0K4xdvYDgvVarhePepyI
p22IpCX6DBBi5xdWRToO9nfYWuLgcCHZQHQ3Qnqq53LFQHN9bzGudJ+JuCDNarSbpn3W7ULtZMoP
67/jUR44NO3K6LzF1XqoZUBzZhRh8+aEYsqd18ftPNrdUQxi50Nbg9MYB9RbRqqbizc4CRy8qSq4
IE5SL+cennhE+LKGhs7C+2htOBfpD61M+r6eagdG2ZNsZjhSclJUJ0NaRti42cTaLktJEtoRBNFA
BQpTmA1SSWqHzrS7HGrpBH8EsVNVuPU3bToDQvarPwwpSY8FCFmjBucxgTEhBzYqn+ZOnFppuCiQ
zyng+vzitoMiaJt0DJDSqABZcmSjHWKYE8KXoepEpyNh9TVj2RykZaZw90tXyCFvuwzE8MOd8Vi5
Mq8sMXQ6U7Pr4KEoDcLRlnfh9TJm8IC2Y70/zXXtiCiv+cH4Am8UAL+BdEBNDfxX+1aPPm4NU+yu
fiiraRl2JOQfXdIpB+nON00e0pxqTzignY5OIIDxch4W12qKQ7yRJT1spX+PbnmZFJkekVcVvUVO
+wbpLeAUd9mOPgt04OaXLnRkg3gMpP1d95/f2+9lBE0mC74C5FSlLOR5jhwm2Brwb0y7UTeEh6Zi
V+dh9du23VOvqxE5ARue6MEuaYN+Xkgcgcn7pYtTsIE+QEPa6M6t5HRK0DX84fw6HNj1Z11OOU6M
a7M+HNpB+9Q7bKBvzYA1Oyjac3YZK0AgYCC7mwfsp1lvGkGveZlVeqTdLkSm0JfWxmjF8XtBHo70
XLALgzvq6CMjz8ng8opL43+eF3JR4/2R3yBDuGDYAI7+3e8wpPRIqCs4lc1EsrWjLBUd4W3DcGno
CieITz2R6j9Gau1dDsGMdpG+SD4ZRLSPc+yVpwkR/Eshnab4d+nRq9DAQKCQwcyGV4EdeKQAOWle
UMLwF6hgw0PEYW9uJwZKewH6R+jhAbTmrWspWRQuTSKzAw0QcS2QvSOIHIGCsp/HfvStnWvVR8Mq
IGlUziMO3fNf/tHtpmYKSlgpwx95Mqrf91PL64/LzNP7PIBiUsgppUMIn3I6ewyRgUcT7inOqw/p
ws1xil32UT3u+qPwgBY7UrZ0k3pqd+3YFBA60CHNB97HBuJWlGSKWjAlXYCjeAtjL+lCy6xcud2D
g6kfYBMBIPD3vBqYeTIO1lwRtJoauu1GUMgTEXcvxD/yQaOuFM8W/gWJfHQ1ohUb13oEIFCS4JPH
yKcO8jLtuTWtyupkDNnUcoj6EeVjmPqxWzLH4YNysAdl5JwX+H/+UNdEwoZoW/gsuZWU11qqG/IM
UVWChjvXjOlJVaa0Qp9w+WdYe+ZagjX3mVDF7hW2HZZrGhyB1BuW/OTr5aU8b89/0VR61rfUNM8x
HHj99XusQJYTp5Xg9y1zsF5Hk5x2ve0y+2Db0jnD3k5gd5NkExv/76lTvDmAr1kvAmocWOOtC8YZ
mKMGRfU0aMhv/GmbMp3MF37ARavqlHzzwCmKhvctOfCjhbO4wN4GJHfoe3kJv5dN99WF6EPh7Rbq
6tIPvObNkJ4KNQb6yAoXtRfjZ2rIQpQifGa44SNNdPGL1u3RzTPP46BKame5S53KHxyeW0fPGWAM
8AhLxJ61S/P1jH2zQquY9SA6QlJ6lQutZsWBXumlMX6/v11MHIXEmG39H07GNUQkA+1DEiSxf4Oy
SS0ZLclNJFzrCPEk65p/nBKeoBur1g/18IOD8LCaVqtHE3Ae+67n5GJQhhsgrbFVMToJ0GamFwTs
Wips2V+qzDMzK1mv/fse+EcyTwGyihw87tqZ4EUYlhNHyw0ApoIeQlsZ8jgAerLcZtB/L3CfnPmq
9v5mcjUnRtLq2g8IrGi0EXtER8DiMpgDKeYVtY4eKg64Lq7WnD7wU1lYaN9jR1znnTsqJWmF8FgB
rZ/92L8CDs3uGXTX41PiTC/DQXr1CYpnbdrubIKpfnrDlhTU1hkTc5HIdrYrfHm3PL1fN2JpgH49
V5Swrs8GFoE5XqYTz5lLM68JG1xf3IfdLV0JHK9ZPRoQItGW2bI8k0217FedJ6C+Y43no4GFX5p4
Qx2rd0LPANPc5ttkOsR7o7cUjcjHvg2//dTQknUOw6s3kdpq/sqwQSd35Uxqt6bvYS/xTxnZE6un
MFDTHaDjRHKsaU1jNyedh7JxwChVSkMi8skYgd4qifXpbwjNXrtUXQ0vhpRUVpm8Qw17XQuZ7fHh
BmIFzyIpITj1r+7pOz7lxJ2+LsbI7ZTp5rRZ/000HQpBVmjPLGT4RZLw8HXuuYkjgodwiYrcsw4L
Yr/ggWtVmsoZmh9l+NOLVNzjt4wqL8sITqSKI6f/yI4c2QtAshCsx4sR5Jk+pXW1i4WpqgayQPrv
/OCXjjLmJNuYfqE85O1IE5cehDqFb6VFEDPChh0Ol4IDnrHlL96q3olbuGRHA71eDxWtJQR0b5sI
/sscbGYkxE/xhvtjmR4vk1E3k+MfbFcCHA3HNckaSoTZXfg0U/bE8R83Fv2ihyiLLb+Zq32P8mT8
hIOoJCy/mKzJBm5lczpCd9GZjJdVn9+dSNuQoYWsGHrBe81o6RPU9QijGBXLTYY20xvKrOkExrCs
HW8xrWdh8Nc0A1T94pEG8sxQ9skvM7HDUrJVTkbExx6d/erYuCSpiIRt+oa0xsqDUmqwxOsQNyeD
eL2wK//12WY/t5gnsPBkdw72tzNV0W3so2mWVVuoUbR4rNs16JUkuSkKEY7V09UxxB3KuaFcMnoX
w+t88Qv7v5YH9ckXyiHZYw6L8wowY9Ag3W4iwzSSMWdlXbyNHa26KVKjBoWmLthiqri+OnDjuc8N
2PLRKX6Ecj6/Zh/3CVgWcje5ekHqOKJnZXzGAzLSohxFMuz9cI0CVXY9u4bvhuo7rTU1pdBY6zDU
u49Gb7sRT0LGDHqPmtoXwGTIWXNZymxzsgs3c+G2JePj9Xmw0j9FvwEMa5OJoMSbbNWYtI2B+xpj
AeG5sdysZouPlGbt60ghotX4lx3q3viqxBb8D6AfrIftcQz47x5a0ICRTztIwEcOwN3Bev2jaoyC
dPJUuEumLZVq0FIV9FGzT0HtpfHje8QDorkWOXV5QbGMrqtSZSIfvePsoO/3ZY0ZrwNUKqGISbeR
30l3nSiz4G88uulzI0QarqXaBphcdVzkiINeI5hnYD33zEWlICEQ2DsMDodfKBCNfqFEe3kuJq6y
8CLxl+xyStpoaWhb+kBHOfZjxUh6m3M1VMDQgxkKiM00DFX872zmCadrB5HjIOejdmSmcfNL417n
yTV7A67M4DLgseP2YKKUYVSortw87xiSI/fTHxJ8qFlrI2BmK7UT73cDPvZZDjBDV1rx5o+hiI32
G0EZeyT+2tLb4Q+ETeRQFbzGugLw94VzCPSwu28akNySrxBYSsEful3kQcBre1QEOfJDYhQ/9X2F
mfe2qzW680LrmcB1boYs0zKK/8xMFqToJbGT+XAT+dE4pLdwpjtrmRCuZiWIWhmDpCxus/2AddBd
KOcjQO1RsSsWS0M3smefPNsa1V3gIM7qmBlChq+2sXZhe3a5+vWoZFVyYmTU/4hm7MDTNDhCNUMd
eSXyfQo6wHdBygJfL7GPvW+XFSwgNNfte5mwrMNTm9JupQHXyUZKyj1r+pVszBVKhTvZZz9hqnfT
gaYk8DUE2sNDyMW1rfhz2VrpJ9asTye7YmnBHFPh7qjKX8hbAaXFZDtMrs6fo26CkcAPD7qq6Eh4
L2pklAcdHsPXoyP5+huQzRnm924nSF2GR65H4hosIqMwpJwcdSLro6ovzZpW5K6fRLxM5iQh7qN9
YACCthfKTKhbXo6dPl7dDIrteTUsUi3fi4AW6GBn/hiDzlJRMELsMOgcz6n/L0Unn3dGqGkW6V8P
7h5JqJ7PNjlOkUJoKRj2BkVrZOkpIuBkgtQHhGbINUvunAUsU5G8rfpkv+z00o+xXpPP1zTIIpyk
5bSGkcySbgJpBNM1+5OhaREkXEZ1TJMmeMTKPPHjMD4w3AL3NULQ3wDEgQgEWRVlYAiSUoZUkNwk
paCOJ+x2lzpZ/LuADEJnzw88A9WZCuIFp1qiHjIguyubyReckBfD+8p51FKnnzTo7APvymstqPa4
dwtng7f7DLfN8fYDIoZ7Mrfs8pHQTox4cw7VxJMP0SnQ0NwP0CjbmZ+2Mhy2gsywNV9aJ4iopFLs
zhdviGCXmb0RH+70r4VNDR+WJCZCGiVP0rDCTpdimXsjnq5OJJRZfGXGDYuxVb/TMr76x5I/YJK1
12jL/tmbclbRO/+qDRfSm4EmYH4/2hBwvhPKkRAYRRd1P5i7JE6JzvGZY5tC9C+E1xG6GX/rdPU9
Sm2WM/paV4tVTDwF/BW74tP9iKLwG80tERvSpNyQ2rwhDF7GC3a+YUtdgHFUgr6cY2y18UDpTxBd
ASIUNtBy2P3ozboykyn8roYRT39G4Lwn1x5VygNm0kJYWeBdvPDbuYq/hWrWImfe+jkZlXY0p7c3
TbM+Vsr+1d6ttuFmtt34y+vGWRA5GHQQjdAX/KWTTrEO0esf+aMioNFEbzhWiuEKsbumM5jsf9dG
woT9YLPjDhe1aVfhr5udHg5YO4O3UAN/A9Dmo67pFdxS0Q8e8uN7PJOKxu+uY/Ct7fydcIdTRFX8
gCrlBHrE6VNl8ngG3QnB+bEqrMf1GgYcqbE2Kaj+gA8kYgtPU6vBex3gY4gVqrUcIxcS4xrLikp+
sHtV6x7iFA3jjnbGWXPDbMI95dhsFMlZMvFFVKMCQ4PPD9kjuOYmzgkk8H4AbK7NcJh642wlrvbJ
9gwCoNeLyIWJNkHAiFpb9Wlyg4FWQKgkdntbf0bGmMdLQJ8Fpj+IlfPdEk0iSbfYGA9BkwQLBxyD
+4Si98O7uD05awfxu0tFErJUM1Azb7vtxXKbdtcpfdBZKD6ZlDjTSnqiZPcRWLajg0sNa5Jt4ICG
Vd5XfSGQGpAacxbyB7+hVl3zKv+ffvi4smDvQhAQfMLTN/qXd7y8wSN1nl9i62A5Y13vST1nwXlr
hfxxg4WnTJSmPkvhauZRZFGMGdmlawjauVcYhMyc+pvYdJeYRtd0XYZO9hFXvU82c9x5LXFBy/xC
mBgc+AJnHfVTu2/WeMfPTWa9rAEqKtSHQiWaTNjw0VFGgY+yJoaXIYG9LGBs3R3PxNpOcHQCl4o4
qSlVJq1YmZ9b7myqifU8SjcR9QxPZYf7A0uahKpz+P1EabqltJNEcEdY2oJkC8ey5xOcNbMMks0p
2LVzHtGphDYuYrPpcrh0OWxr+AAxdOsxoCY8efemcnMrBIZai1/TU2u9Y4/O4VstMGFPmBQfzLTn
RShdSCvbjEydeKTUT0RtAkGe01z+npsZTfPnUKA1DOoRpMlvE6mc/gEjTAxtxF0j/VrwPM05k15C
9NZq+qtc+a9CXENNILmEhebLbI6Or+rXEabyNScOsHSZovlL+C3OjQhHiPiLUebCCGWFu4wXXeFz
wx+NwbmWjAF1tYe/NwaEcqmZcWRl1erkh8Nc9dtkopBgYVWoOKtE+epyxEHv/MP6AYHXRUmfn81g
9uwPKjPZgwql9L84uPyJDtFY9EQJihKM0REJXFPQo/TxxdFceMuSnjitc/eyyblAtX2LJ/14+GDA
F518F24ahLzLry3wQ7d67u9bTKbIs167My4B70SMWT6fpR48RNnZJibqpawPuzXJ4W1B4SoAi4h4
MtOMm8bg04eO6tlXvx+7R12qS2zYpwPNuLjIMR0zVmq9ef0nL5BA3Bo5Ez4P7mZG4G34gTJyK878
Y1s9wQqS9lxxYB05e9HAN6th2IihmHgZOu1zRPbbwpXLrspPtE5gKbSXS8umeHj0ONF/bS69PFJ/
3KjAeTMnBaYlEFCIJ8DYP3HwmnR00uJg/Gz67R68q2mjskEv16XferScDS9KeFclPWv13T96wmoR
eOw+H8M7dWDOAVMTTX/XY6fF7CgEczJZhs7l3dEveL7sBvmgIdDBpvqigTAJAgPEHh3p9llN3xxR
I+gv391mCdZR1apzDIQ2yINDlo1Vv4194Bukm6glXeyEATz6gYMOqWPHTrOB36qtOEPf9B9lXXVG
caDqAeXkgj88VZvFBYLRPBmAPX3fSVN5oUkoE1IsXdgfc+mIGsltG2CKe8uRW4CALkW6V/YM++t3
knP9JkLGpJmelgiedodYAJMU7MOO2B0+P6+kY0VxUMaXb8zsHaIrUDt8kO6K8T0xfT/dwF5MP5VM
XRF/ff1TujwPlt64EXhItzGeAbL4f6DxgYCCIqTn7dctMqqqoaRH0CBw8oWUZaCssy6naqBIX2gI
Vh+FUQAJ9wIlTAb7T1Iuf6ciuFEmMKDH0w0exY5I2fExLUkxXLqEr5Xng638PXyXfYMlcXUwCFld
ImosWB6P20FU2SGmjo5AIVRhKavcQETQtoZQvmtaCr/JnvWS7zHlMZ1d/OvdGb5AEyhu+Xa0hQF9
TatcIDe3nVhTV77Yo4Sixty2+9QMA7qW9aiyNpKca2gRpXU5WlZcE2U4X7Zi1UuI9rR4S6chrrGJ
iHFIcN2ffi2wKmNNH0sQReOClQSescVTCd6YVmOQW3KVKftJJ/IaatePaHjhb+IoOJNcv5tuwttI
uPwH68kxQ6qzGONdNrNw65IjbVAhEmNWAgyuHKJ5nr92y/sgHLQX/HZMRXCVTng8p8KxW3T6FTRf
gKYJc2gbfHDpcfm1KmUnFSrtytjicSACLI969GT6YZmH8UiAye7lTRmTObVqctguAGp+wozoNzdD
EMvo9gfS6ag0daKJfcdQKJKfntArToDzGx5hrMDY2LssTdhEDaQsJ7FJ/PXXBMY7WAV+sEPBiacz
A+FUckhCGRCzNjqwhIBd9Mu6NgQRmgZsxaojNfTvimkseNe2JnICuofrNsNMsOBi1Kyh/YAjniNz
iJNvHMsW9rRq76s4Zb+FEVhGVLNLqbCQHQX8mBKfeOJndeABw+tdUIoAVIoQadraw9ot5XVQKBfB
wvfpvLYfHHU4/EpRnRiZGtCpSauHCkyA32HIzUEU/+j+26U/KhkxTe7DDE71z3U7XxaYg2rN0kcR
/Xpip2IHq9LmHVyK4z91n8CTNpAdLCMdUTpw/V/DaNGhyT0M5qlgPNyyyJqfDQRVYeNF4Y/lXwu6
OcYKrHYCmGTFAO2A+bbW02YZXBYjOqvthFQ7xFhoOCiSFPKsmhvEFfwKFHEXxZSUnQwWDJ9oO5nq
NWtdXDdZ5Ylghe+GRA1GKoMt9ZWbDU2ZJK3h2kBmTjT3XQXxTwtaZnjrPLjD8eN6qrjd/eSgTKwd
5Adtz72NxAwqj5pJvVPlbktwHyOAAAKW7wKFJIS9t52iTYF63/6hbTrog7PcYhqE5zhRdmmGM+hc
xtjjwaLb/ExoflFe2vlSSG7fVGsoSAEdUsQOAdQVbbIla0y7HqUHEn0lMlnhX+4YQrT2gMnZEDLx
ilT+n96leyNW3mjmvwI8oAAnN1SSHed1Mm9NN/8QJ6NDg+eFDYInL86MyKW/bu7SRppFMZMm5W9c
GpJ+5TGz20OsdzLNiBzMAQrrn8DTD3XojOuhrLmpfLSoniptPORPIy74sZ45lgLd/jxaSfnQNFKi
IfDEDWmfTRUqD7Np3UkLv3XUbSDLmw4v9+I7R1BCdmLfD7We8jercp9xqBspCZxP7rHfGarohJU8
H27svSpwQkxUfqA0zXh3NyDkEXc9llPPn8BreDbxdT/q3QT2NOoCiMK2eH1ErNxDvfQHRyIVXDH1
ZiXd8XzmDouYP449TM5sNZIlUdVYsF7ddbcIrcPKA7Nnq+A/AKak99YcQJ/CETbDGFT58JWFg0v7
v0iD68u73fTOrbgIXUE3t6bfcDwPSQvfNCJq1sThXNpcinKoGApzzxRrEddzD51jjMY1V8a0xidh
khp4n7ZREx0duKiLW5BzxJpO5mw9fd9DwiiapKXxPFRz1dXBJSJw0rPB+DVv9L+EEmOdljJOmC/R
9vGZy4nlXtnMMrktqByZKE+iSjC5RE2VXyjJw4P82kBoRc+pD3+rzIBC1gP4KmRl2u340wgqbBos
adLzXN120duYrIPKl49ef1kcXPEsDEDqO6l4f4H+50wV9kDjvVkXm6emliW37hhOADCm0Tje0vFB
W2whUCh3rXQ3QjNVT5D4q0FOOTEHpRXc/ePrkRrphVSC5TF0hBQmquirwhxkSKpFqSZlo0EzfdIc
HCY+wcn7n6A2c59kjZphhBFMulcwlwdmhE+RVo02weAaYP+nwusLJrm+zU71jBRN7Rn1PJcKExS6
pDWhW9Vu9rhue4YJpEWNksnrgNSR7zdhlO0ei7eAOdN6QY2ChMEPZWMJ/CROTZ06s6/c+srU+K5j
EnfDh0NhueqkDNauixfSUEkzg4BKJpgXYmoz1BeJ+Vbn9mR/syKUkjXhIshx3DNuLgRmEBi/EPCG
2BQxCprlz3SGvc9I3wR9NLXfCj4WLwShxNE1WzVxNlZ1uSVjaupMi8YU7CZth13PaKIKVcRMkzG8
O04dGEcGA/Ic3UunyJBx0jWtUgbMiPTVfv6f/z7UyRzIogs/lj2kfvuJc2938IuFcTYAyHrfeYuy
D2Nh4lbMU8PMk1c+FMJX1eMpf5VtP0hHgftCFkYS3o79eEPi0j+JX5cBEu4+CQgCd1NT1ur503X/
n9qI5NtPb8FjIX9YrJgOkZzadYPrDPqXAayVHvrV6C34Deoj7UeBz1Op4SGDqB/ZCxhHgfmwL25u
10FNfpdf9m6mKSWtd8QO8uzGV26+9Xcyap9FwutF1NTuRHx1+dCb6H2oVm59kgyKJvh4idyqIJFy
ZU8cPcu4JeZKgFK81tWRz2zX4XtZdXju/4nUjnNPWWyTGC4TveA98nBNJnegau9WuNntT/q7EZ33
yLPsh1b4NFLs91t8uXo6IdeOK94w9djnURMUMM0QcJPwSr/YHNoisK/3zGY/oVCsaXLHGUHyg5a0
sFJN1LFS4EbfGYCJhMm0juLbSB1VrCl+86w0qLee0pvyYWh+juHcve9zenZXAPoQHM9XVFddG/Ez
ZRouIpTCQqmkgcUROlVSYUEmG17pe82g+ufkIDEBhCbaHllPnW8huI0+buHNVSIC1mb+EfzzUZ1d
hDVVu+mIUOwMcJixJa72TjPflSNrfhg05V/G0rjAO7JuMAtQLWSzWYHVe82kXJsfLYNTwAJpFwez
k5+CPG8jw++snUzipVC6H4WYtYE3xl7W7H4KdQEJh2ia1mU1Nxir3VymqIpO6Xsa8AdeC+hvzW0Q
tUmyX2pGi7jCREDyVwUHqsn7o+uonuOBij/VALDFviZ6n6fMHG1ESl4n6dX/Grs8yQNBEgsTfC1G
INEJDdV5G0K9Ddc4EpwlJVIsmJ4HN8C00o4nQC/iI9MhtawA0wf24yKd9JYgnTEejeNvt2jyuj53
hZayUIPDyfW32AUmR0VksMIn+ZbQMOkSbXgWRrGPoiZiwyVWj1HJg+rq2T6uKaN3uUQzBDfc5nni
2XA4CG325YjdRaV199MS5FXjf80pQx7NORGxc7Xl4HpaSfUz+z12E08p4ro0LwJISKtTte/jbeM2
y1RD2o4vKWW6ZIcnHhMaPq7g5RRZ/6HaU9T9cu088Er4uJtwbtNv+1XvOJBHD1M43mPQEFPZlD5B
ftwN8pcWZb7dNUfbuUCaGNyyhrO9TRBjaXpfFlQMilQzTWwdA0wvHoRbOcyQ2w0+TCJkqydeZQjB
VLrc5lBMpHpLyP0dApbfnbRxcwxS0ZTv2BdJtEZbzYSiveky0K+4AQuU98BKqgAi2uCGfiEyd9MZ
jZbd07Ymn4aSJ2sNKnjiIlS0247hRcKutPwGX1fBK5v1JjlgsvLxAP1sV48wIO2LUjnTPyQ1LOpk
mkdumF7uNnP2tTFLqP4/A6X/drmUvf0Ij6f3ErUHe9UimrNJXd+DVsg6TF9ilhlU2URhfwcovCOk
9JR+FTwJwzp1SfS5X/VMpgkqEGUnJOJZhw/Afdp8EuBadplME0FlBBOAA/tlSz560J/kjWtUk0a7
5P6R7X7pF3bWT/KB/HfQvKkmZDB8oQqB2fRXW0VCLeR/AjANVBrau2QCfxAxEtMgarVw4lI5egEm
/auTHnSiTwtvkRHkzI6pWwCVi8aIJ0KdNhARVYQJjdxw009hNmcnf8s6kK5GQimmge4SOjqyNbYw
h0+nMx5hdrdOEZvCWNMWeh4TaeQ2ikTwwpS5YH41NzvjjYQtMkeAPZ7HVfx66QxN3Iavlfw4hkHx
oUX8rO7mR4x8tMp0GwjVeqWaarl13YUGNiZprss6OrdUzyFyV11rmQdSjgz1X35Yl7bG4ZA0PI/z
MNkZ+IreZvVteZugq+gwuJQ86uTqrKFg1vd5kovHXKVVE0PxXR7fbHmb6Hb6g5gnigcF9brdDZNe
DyG7MknQUfP2LpfBQnI6c6qXYeLAyjpssUKJ7Ofg06C+c36x+Y1thPmPycAcKu6JIVLT8d/xdQpV
9Yv3NxWdurORt2PnlyjD/ggMZGI6UBWiMGw+VsltsgSWIQZOtfO0dfbA9cr0N+dKUuRmFmrU/TgW
51GxBx6y3c1qg6ok/HInzoU2i4T+SCTWkokXiB+Ukw8U4ryNXApLTo9o25L5mumDGJOjyMe5BLbu
hpCgx+kGodvge3dC3Hp04qEQkNxfbor2rIwTRmVYtBj8OZ9q/YwbQec2eg767dCHJtrAcjQzVvDR
HRApmQ6hh6TA4GRH3CQGzvmbDWUNXgM33qZeOGFeVcJ3DHqQsbvSg9vQAU9vAZcm0CNjasixMryT
a7mk+kE8vU8mwXAaSeZJOQI+HXToOrr2TzZdgQTGflnMC8/G0pNWStFSvhPHeEYQn893vxA7lQIa
hhYlC0BkOOmO8bloMjzQDIXKYtVcvPkxKejCXiM08bI8E7k45vUpPKVdFTmpkGMwrkzOsd/UwR2d
ES0AxeNSgF0IkTAP4xt7BzirqFFwpIb4kEc6leFOKy6Rjv/+ZwjaI3dqKS3kSICz9J/4e0zYgMCH
cr9bB++ctilh8eDynzRC/FdA7Y/YID0mqt0HbqEEuCLkYfu0Wnk9yN1P86JW9fqhomgcAdSnTFFC
oqyy4xmws5SWR2JD2DWyvUKuO2u83pWZola7XAylM1XUBqtzA4u78rSfu6asswSKeJj90BxJtVBC
/Jk4xsBfA/SabryTpcWUcsk2Vx8BiPOemj96btC4C8HAKzF+5JWzSL4vzObmIclJ6hltKSoaqBF2
UqMCOXk1eXHzgCLHtcza72eTL9dWQw+OaM15Fm5s1B0g0BB8nU/Jhq/s2eXf1tyF5kzc45/YGSKM
1n8g5a8decfz1C6ijJBn7a87+edMER4SdRQNIyVJLtSl762Dt8cee8oYLslLsVVk/a96ayX51xzZ
dz0BwNRyV/RYq3B1vT2aLe3/GDFn/NSYYAkHt0ugs9dQZ30Ue5sIImQn4eMvCMSV8yy7fEjNMq+8
tH0S5RB9eWmBmFuFLYwVbIGTf1G/UeWP3QT2apqfGPnKxu99uMqw9LBP1OrJtixnvHuh4ptm9asv
Xm936G/21c5Sfe2e7clVOPE5RXz7+kS+EKPeuke7oB9JfBxp48aI7EhVPaNkVPK33OGYhoa9WcZK
+QoBv4UfFBvFpcnjGnBUIKlKgABn7QHtLvGagRruy5/I6QLNgv6c9G7FCM9OCkkWRG7eQdnUJigh
yM3p9IRcX05x/hJzCJ0zqK7u1C3a+/3pcz41U4XO5whq6tbw4wVKxE/bwKvyyRvTjh/wqpEXBMk2
zNWDDATeQKoXMS69PsQzN/uP2Ty8tmF/0ozgvWcKmPsByHxUbxTzhB2odSti71JlOCrN453EJqx/
jwmWvysITQRNTuhMSn/BPj5xTCz5V9S5UGPK8oxCqJnuNrcr5bVdpH5h/MIEbyg0oAivAPH8fN+f
RiOvRUM8ijTSehoMJ0DmQK7GfbnEH5h71Hh8WsrubPcp3Zks0prt9xxRnWT7TmfUdYzBXKFDiKEG
60a61K3Gw/4FU+F5yFuoc3GhrsG/OxmSU72QseNNApsZ34uEnWr0fXsHLKfoe9CVM/jbh+ctZXCN
kvfgxesbKJFSj72eSgzPVZeuesaRJ2DMbf/dmGwOZbDD57gxfHP/vzAN0gHc9TW0q32/dPOTVh5m
3ywmFjOcyPAdNFr+bXef2mU/3hB8/4C/1olLR4jXYaXFF3460qVphzhEeS3DB8aVYlikNH9dGU/4
wubJxC4nUIljzFNy/ViOcRrmJdy7gVIwaOCTCMbKoSfARH3PtA8T2mdZ3+m6St2SnpmxV7A1rOwD
aUd3oRob/F0P/HxZPRz+Usb7/rfQvE+E5BOXvMvqsZNbeuKxP4TsPJt98TUTqDvqp+NgJYYirn8s
fK+j18Ioi3PACxFAFADA4EncunezpaE6Nn8QOZCoXWp+tR9yo1x8lrcS/GyyZSj7sje7gfBEtWSW
ktDoqWultGJUorBASLhFxTWJzHNMaXd8EkZ43+Ig0+dOYYkeDuw4BfZRd0NlOUj1A7Yi08fkbHOn
DGlQWO9Yp2QVtiRKMu8JX62HWqdDkKKImLv5hd4fQtuPY1HW2cOU6YNKFTsv8j5b9eU2jLNPcSN7
oAGmuuGKJjeJRRJmtIbeIWHMqnLETIZT81v36hPb9N7xwc8MqahIvxyRxN8l+feEijt5AavO1rIp
v9gMTKFGuMfn2Ft68aueU7NMwWqnT9PpJ3QkLYWJsa2Y5S2zlxuyXSPaVaP19DWfT0seoSim4Cic
PhDmex1xkdRh1KnPUs9qbJKJ4SaX1YgiIZuG01UOsbX23vXODAWlEd5jeddLOvriWyR3B+Oio8RX
RG78jbCYXRkI6KjaSodeUvoL3krjvVqC72jGVscgvQF4iHf5Mb18FYqxwj3C8TbIqEZbs/dQ2buZ
vWtpTiS24DCgMJCb/hYVFnhEPwVyGVFkE8Dfo8wFgx4TG9o5ZyxcheBKZ3ietJIxQGOwTW1dI3iT
NKx/OVgkjkTxWucFkIoyisueg5mQ3HiNg3CpKj+bnLnxAiCRZKivXI2qUhrADGzQUYWS/jXb2g6B
tUY3J+rVI0nCb0ClN+aOEpkbXA3YBVdz1ORaHAoMJPDTtCLfkKtGPYOXr8uqFzTiZMFFyAqYTsQv
i4sqBZALWT5IDY1H52PoCNVdtfN307N+KsoCgqNyz3JhXQ8SKpRYxl0EMBFxjbNPH/nWDoHLsfnI
+fYTrVI3ZxQvcbCGNv5Y64LmnCXN8JR0FcbsJPni8QRTl7YZlSEd0t9dNqSAd14uuTLJsZzc/GGW
rn4Z3xUmzT3SObrtdc9RRwCHuUQJollIVmxa19BBcC7gwvX3id3rdwbi9pAkNTsccnMBvaegWNFk
VrGghRARoHEYX2tm1Z8zHpILgfFGhGBUpEjhGXr+65wgwqJJOZXDvt6gUyqM457g+ZAB0gdZPApL
e/IG4ONDynGMHF800N6RwW5nq/Cvc2DEsYZOOLVKABOmvi83U8WpmpPWJibIxdlrsNjvyXArno5Y
bkugoGmYouGCj1ZS/uVNRhrD2k5B5IfNm7enNh//jIZcVCE5mN9VQ7KXhmFaihH4bYpx8UqG/pyu
c0YK2T9S/LPTkqlwNNpSpE/lD7ri0ua9nIsHeYdujW+t45WT7MHgKs90Cq13S8KGWlVKTSPc1yqW
jVnowUiek/FC+KehJbHnaaR0Orn+mINqmlhwOuOO80g8yGBfuwvSvq2PpBN36RDlOX9ahXsGfd+k
z5goliitJ79wZS4Gcr2QWa+KsbH4lipeA1MrU6XOVbpg6uCKXaJhKr09k5ja4Kz2NufPpvTgWQuq
sRCWleuXDJdpKZHMZk4txMaRiGdY/k8PjDKRSoMbe365nbBoePgFkzBC/iPdGQA4fy0WVlcZ8H/r
K9ZFUuyJ4hoKlN3wFMRYlcSWs/HtuqbpHIOhxwuow0S9JHeo1Dr9TWo17nUc3mSkXnUWdgWditk8
LSqqB3VPnY+LxyiTG/xdBnTX6Btvy17BXKru0hLMwvuB3j17jmsT9KQKdPo4XFcmr8EqD81wh8fh
rOyyYPctMFsClQg2ZPbIZyOfSWo+XJzBliGgWx4X0dWa+fpk+3G5Z9r19Isx5S7IEEFS4fJPcFvu
WiVTyFPxj75IriJ1xnjo4eMQo6Sv/xn22ta2aY3GKrRt+euLycs+Qh4qJ6uxtJFsi1gj748kZSIY
TN9CFIgFoI3USA00YmMG/NkPH9d4LGwunRZYfxfuvGauve2nDr6w4/iDCLDfh4My38TC2HHlePlP
sdZMUGVtJ5Ai+r05N3NDVRYPE8WTwtmQs3j1rd9AD0AcHk77zJw4eTcQYYdy1RmLyMLLL3nTDlrd
JVK6WENzlpDlC3PezNqLkI/l72wehUFyPh5V0uDPOVHN+YPEKHDh01ub+jrabQg7mf3wZMH4T147
BZP3F60EuuTXNaunuK5oZamuU1j7nY9EtPAZGpI06xmES+wREso1dN7fXQXb1KU6WopCiQrfDgp3
yjlDfwL6RWLCjcEJBIItS/rbXm5BIqY/6Fybq2lUfFHeuQ4ECoF5sG3dww4b3dw7YngpWSSpC395
nWm4BjRIfhvjG/WnB3x68/1ykknTB2Q1vS6l5Jucxr3PJoIpId1EuqzEQr6UFOGYkvpeRqAC6WHZ
aGzHUWPhAsaUxtL5ygAdg8Wgm4p9W/tC6f6vMOGytxJ4N7rpFWqnoeKirCjZ93ulEcuaES/sRBwe
Q9RnlWovIuX+fy2frWcHlZ9LN8rd/3OYVic+S/CZq9QjuUo9FLwGTSQk9E5FKZym26lrBK9ywzvK
/RBnhXZIuBP2JoxFMdlOTJiDpxmD4zQDSk5YWIc3+HZyvpRID44UZZqn6rXhDeC/rQnnEm4Nn1gL
ZltgjT7zf0NMMGrdkMX4XUYGNoPgXt0FvSnQnuVJIcdpF3RLb4aiVZ/ppjgWpdYBu1gON7uFv72G
nlSgonQ1kcde768x76h4nmr0YwtauTr6dMD3PuzaYoStvHv2FH5Gt5Nzt02Ux9AwjWnoepHATtCn
1ZH5qcAgfSvtCWuQozlQOlqj4qxAGTNy0XM69+gol/PRmTCWRImXxAgaBkskjzKZELICNfP/oUZJ
AQfgR8zzn5WpvTJWWudCSHG/NOgIL2phHKVoy2dDYhuKTjWI3c8sTpSZQTVgZNVGZcYl8HyxcfHJ
5EDHfElF7yYlYAFDzJeUOHxYAbD3BIxmKpYzlKIruJazfSsTB8fiyCRumiypuxvw6GBguu1qOmQy
nW8nkavXJGekcqrBkZaJKRhGLnpE7t9Ep19yKetGuEWwHD1NGRE7jHVN/LS5p1GhBi0iRc6HuhOB
yNYqqFVXCS10aPPA8hcT3vcTaQRFkvk7SVvZLzqyEwuDy8D+SY9aWJdVou7auyWi3hKVlF1eFfve
Qf81fLUIEWEDZo3geDs/DgVEIKc9TmbRW2cqUscbD37SlkdHUWarZYEisgubkggo4Ypm7ZP/ubrv
/piGNlMgkPkirWh2Y/cX8kP4pJPkwyi4wTLX+7uXAm5j/KVrPCtocSlc4s2QpRvsE5iv1JcF4Bql
wTIUcxqoBSZXV6+6KbDCHxvOXOnla6VT5Bg6H1fSMsTmKdLcn5dolXGMzzWMcmigGcUNqTtulXMH
rnnr2r/JBkAqtfYGxt6xavSHWdTIYva6msozBQWBkR6dHSVXs46d8aATesiodW4wIpLTffRo705R
pA4kKzIsPLv7nPI73wgs609kPmkz+z8W8J0ncsxvRoPDOF9XHWzBlnGjMeHr5eNO3NUka7DfEZzp
tf9Brp+l4vrZhBKApoi247/+XE2Fe40M70wnVHB9kV3Kp90YFszfeXo/WhfsBLRHrRdlyGGDMs7t
1bLq8RgpK/8S7deBe0ZgDHNKKqy/dV2n9pZWyid9lB/Fdep62ojoCLTVzzwLnHi8pqSLo8B5VUG8
CYEfvhB51ptQjtQjRIAd62HcxPB42nHBCkjoiV6JioxAtqGspvU97tRfIeVdJofrnYgWUHKX6xiP
l2K33STRG+vpPPq1uCB79V+JqmlEDxjFHp3h0/6I1Nf0P8rmJlW6YYW4fhRPFVlu3lGr3VZD527x
rIkawCYJMk+qSx1+zObaHHuJK+L/0V3ryjaELf98EPKKQhnBve4wjYEh46Dlv2q7N2p8NURBRucL
yXlgarNUt8u9EzlsRXNEYb6S0Kk5Co+Z4sKs1aGCE5TIelaHQTfEYlntpuSTzA4q6GFqhU7irDAy
1HHZzhklzCY73MaIhp6MMoyF/B9Gm8ia/Taj3a5vsjV673R5aYAQ3Nql25XgWwkS7TKfMH+khPSt
9H8fBz9Wb+Kb2tdrtijLVIda+Oy7WPtRqr77oONUsgEfOOmzBaCk5TXJNwYht3Xqo6+XgHkxBDk7
jTdSwmC+4dVzplrJNnITGFE5SY5XaASKyATzVxosRIlBMRap0IbIwK16JlKSB+3VKaKyuc+cUHf/
hTBKcvld6IlERO+Bgjpx2N/outvN4fdDR1z2JTV/k2FYhKUqIXr+vzUOwa7d7Y8RoYn+0ckB7ZGh
eEoc9VRm2kHUuDfaX7zV8UCYGweOrfrPDkn4cpfgJl8sjFY5eH5iPue7bGXBSX99mAd7FnTpNeUO
VUPwh9ex61N+66OQiVoxI6OLMKCxaiJ0//I0lSPcHO2UBUX/xSPXaoXSA2mv0dDQHhsgnrom3Iut
jPgneaTPgdDf0Rwduw0wDlGVwbmxRwHTI0hz9WMRu5Z2mmB+zy1TFFxkUxTr335MQZNglziJu30f
J6VTWrnbMYjmpIFsapjnOANf+1yPITBA7+VQOwf3PXY07min/oZD5e95UxjQ5765gWNo7knRiLTZ
k/EsgtuKxDPwZ9aForp7QZPXTr7v+dDUTG2nxP48kB0eELMCN+HuVZgIHaiC7H2gG7V/BtvBVAFE
ZWZ+xJ5aNsqJCjBASWvIdbE7q1Xdt5+R/7FKRQ5fBA0EfrwnT6RmOt+hE4JDNk+DT+jZNgE1YuzZ
BZgMfstld6RSuLd7hzLwwky/rqxfHN8KO9lspcFK3XmCPqXTc61395G1x1tOvDzTlSStCJWb27GT
NF5wtaaLRzDW9KHFbdGNiielFVkYKVhVneIhoOX1K+NYzZa1tWbc/3cXWaR0zLKI+DBPWVUNv15E
JI3IzHuMU8/1PE1s/DrOYHLdfxsBf7pUS3/V16ALCqTU4m92BwR65Z5Ug3W+aFKYQ+dLRZCrWnJ/
afx9Tq8yC0drEbOOJijnx3KSSPuUQBVOmXbPZc5ikYW/mqdI5a5wPEPzL+UZVhWFFuFy02FT3V+Y
HDosTfu2IYRSgGHoFe1BCSDroCsMUSVNPJmFk4xs4kKoeSOSAfg5ZTU7IrI9v4SiBMAdB6/6kJmo
NCNcPQABwm69egkQ27sdSRRcDyFExDPkGkQUj9lCQ4MucH6Yev1LY8rHoZsyiYd/2lPsLqSrV/SV
VO8D9RcRoYRPLUKex/6hBOF4oPBvzga3XOL3ynW1qEVubmlPU1vdH7jAQIChvUVWnRF9W1sHzxxi
0AF+2VfJ7PLW8p+cetfhKCybXcvp+ig8LB8wfRQb7zdHRHL7GWbKnsZTyp0tJItnDqP1K3NwHzkk
y7BmvNBIAx6IRESL0xu3DAr5AtLoQ9Ke0RpngmDK+cXQ2BFHAZOaWnbRJsWwG4XMxgxXoxMohWvl
DAXJGJfebueUEncQ5coQkI9oUMkTq29E1kFyz05NPvdp0+WC0cl8cTXzA7XdLENsSsg2dlaVwsIV
pnliWl1GEAYf+I1gSta4Lwp3n/hwl07XpzacsF5hlYaQZA6qIEcqmla2DjK7Hjp6M0w+IHHfDUHJ
BFs7fkEfs9GqspQUH6W6sOBrCKsTSDDMJ5Dx6c7PLIMCWS8ZjNYVUdU2HzVCgYjeoU2FmlXp+yE0
q5EGFWyly1cgHZ1ZGStXMGo9uFk4RbhMuZPQNxxgj9UAPLQ9IaQMQhyNgNZKsKPd93sJwczPUUfb
x7pvAs/AZ5IhZwMFtaeo73PoABd0/9cTDQsT77jqmIlPiL1yNULKWHO/CtrrdJN9eOsKmLOwM+RM
deGrlZqNgAM2dkkSkykYGl5PQDzJ06fTnL4C7yCE+ANI9oHxHV2tbLl1z5RA7Neqaie2Y7Ozambw
VVUdCt/RNZIyM1DfZ+y/ug1kR8Rne2CsLiOSGxfh6t26YQi9eYBW4gbEF35iXHTE+79HR2sqsT/A
se34Dr8Jc/gqSdlniICBVQh9klCG+y8oZY5/eHF9LbOxdWSOme28gUbgtm0oyU9NIQMM4CDg8Xo0
fSBxMjjgWUx39Q0d/jueSRivzWJJif3hhO1aVMW0Wa/e5HLYE8P6tXvfh0xhOoiF9mfVZ67OGMGu
CtJpfhOX+CznUBSkyPH2jZXrh73eMp2THFo70TnnhPm3DAQm3eYL39+KAyRRMy69S2EnvADwnak/
sqlVmWoGMSSabbsoRNQIs3+JE/YjdtAv5TgWkvNi5qaym0gR+ZK4a5jhFS4GH0+kBvk1xAWShYC2
Y9y6lG43n8fwnoaNhGOoJXrO6tHgEOHyLL+n2I+/XVLmLQJwHpYv7o+IZjQlmoakcgqVq58OlP9q
edgR0td/4JblsCOjVvBHqT87VEp6QeN/WvYLkJC1onXXQzSyhoZBB78hva92qnKrXvZ4DD7Ok9Ba
/60mlotOY2WBcPPV9vu76xWtFVokx50jRGJg2Tu/jqkmsRMowF/5CnIyXQj3vJ2LtGZ66z2mQU3K
f3OXX1XJRI9Fr4dJs3NR/fMh7Tm3f2DoF77X8gVgBQaL1bOwOM1ozPFctN7ItQpJ80DckUhfXgY3
b4FYX3iKWxg99Vu7XjxtmhHI6KzSEAaUT1DjqfuVcw2/aUr6pnkMgsjS8NdhH1r+0ciNxVzsuT2A
iK4ct3RGefF8bDgNIdxGhgVU9fl9evbmrIP26/1l6ipE537vfhaDMTRtSvmdETZPGMy5+oWVfqsm
83Cegn7J8t1LELhkAxKctM0enls38FSbOVjwIQQm5H2f9rIotUUd92sF38TRU4ga4mZ96xrsTfNZ
9x4YrLFNsWGgrH9Y4MtwSSYOFPheTt2AzbYaC1MYj53zKksa31Is9CAqhaOScAO0sxyt++zGtvyW
TREhaRZB9X+DU6a/LPQi1VNMQxreFXidL5OAg9N0LMvZq3ve08td4chauXFl8FrpNQRG65qaCTyh
8d3HVXn+Hk5XytfmLOP+x7R6I2QnnG49g55z4lC9uHb0uq/U0ahPonyNZQmI1FUTPY7jywfhSswW
OD1XdAL6x5tG9LnUtKbf2jzyQN8puWi9xIcsbfU9Vihb+CBPCQVOASYTn7MkqO4ljlLuLIHfo1/U
KF1nrKqDVcilKcd0Hc/qt+Q6ivvohQjJqVxnI6owG48Ul+lKdf2Sj0ljijELd8aBf5SZvk8psLg6
lCu5ZccADbvUZ/g+y0+LLfpxNlgtAzQ49+5uKTcFa6K7DPd/x/t2UQ4WZoBYrNHfp9Dx7NXR28LZ
1lDXpROd70M4aVV4qxNraRQ1cnmMAD+cYHcBeGTxm1wWnUdmQbTr2MEIaNtK1w/nk7QIS2wPepYy
YI1e2sVpCgEvrSgmZtr7Y77o23sTo9E8iTtFXIyokduNREPE3QQDxqPgpcUx6nAYbwthrechq7tm
WD5oS2RKbD/PtMVzYRFTDDKhXmTItm65iVpzEPpxKkylvHkR3JxP02wa5SkXUNGaxlEy+k3YGYQm
2tsZqAntKNGZGK9nUz9ouPlh9qfH/MFa4icVSFFVIPS/I8XV3Tw5KgwonuUMltw7K02f9mjKuZir
Ce6g+Km/BnjTlGvRSiyR1hF3F9Y0EQIvTYDd8Rg5Ge0iwqxUZNUe9Y6CSGO1WerFewsLF6fAA8+z
A4O99qeM8uQqwh69dGsyBb4yA7OOPHi4jFjizlvVnNNFUH22c8INjMvNs2oZv/7iGuDmJG21Cw0j
I+X58Tc/Ux5vcxJvMY8HAFjr7oECrmkqQepOFk4fa+GiHbff6caXjWKHxmkikXPpe8C+7vTD2IAY
kM7+08kBAO8BkkMbQuXgcnkC7yJtm8orpIATbVzWWEsCAlmaEcv02tSeTaktQIrXmeup21c4HoRA
wunhZc9Y+yox2yTWFoFDu6nUCyUl/G6Nz1nsncXAcX0lnQFsKbGEQmLxMVG8bXgXU+C2dEbcgt0Z
RoiFWgAczM5kIxfp2gpX8AFBtvT2K6I83UPah+Ftenx3ESVAZa9iJoauV5LSFQboV3ne91iP2upu
72JsGMCBnX22Qnef7WHeEniA/cOY6ePALzewSz8eeLXQXJM8dFE8w1EAos5+M/mzd8qrERb8ezvW
GgiKY7yz+QuWylApLBhEkAa4fNOXTTMhQBARIzkug3Xbh23Vk6r6TrDqoCIe6GM+2ed79PGQ2Sx7
jPjxib0n5zgXIcNiWn0wEBMv7x6JVr4xw1DChrvHKqd+XxCsq20PiZccbqMfBJ7WrmR3CknGc6Sq
y7PGdd3vxVNpT2W0UWEtPmGZOXvqohEKcBNwRxjjMldNCwJbdAuHUWrSIcIENsnuDU83lQtw33sA
a9C+fBwZ2SP503OheoUXjIgTMx+8uEQQ9WrdDVqcEPSmJa/nEm5URl64lBz/fAbOQv8H93rxkJPg
ER2XLW+toSlEoUL/klJotdR9pmR5ZzpAhyFzp4+oWBwTlQq4UGoyfUPmfjmqCjAbQUEKhrQtnS1a
s4ERBwzflLIbophfWi25ZkXJuHkpchSfuVVqcdlRFqmVllC5lvJbtRb1+WeSpGFe5toZQg/7LuXe
YZEkj5TInA4rj2429mar/XgplIDnCA+Kzo/bffK2B6vUeqqVl7uudplMJKaby5yceU5toLHA/2Lz
WqIC9uhEOuaWSRaphVkDOI9YPLa5eb0sc//ewNnX1NfEdB9MoNUAXb33VHz3TxkPD1xNVkHWL6t9
5Efq7ciB9wJqL8InrebQPOPsXe57cn2p76JP6eQVlQQdHvUq0VwHet/MQbNWB+lHAXS19mhHzIBH
BFFap/nPUmV9QnzrnVvunEqJlUVVzJhKPSXbpI7ienppyhzM7WUUQRoDSW+VQgYcMMTuJ2wTV2Gb
JTaOfuR7sBMKHRUh/3u3ixJUfdA7cL1o4/qtkI7Dxt8QOFzJzyTo2UI1NjrXTaq+kr00g+1hM+oC
cY/zAAXvrXHD30ZNtG/QsHZfD6rvHW3jghVvAHc3kRs7jb6ZhMVS1PltpuyoQYUOXXoka/bmbh3s
fZzgx7f00CdI2mWOLaZ4g00fgXG4AgqI944OqwAomrAtPfa5xWHs015g6uCL3HSFwirlBpXM85ij
ogQCYbcjjRRfVNc2Yw7Ov+P2fq2ReKpHbnhs1IDum2PjPjUMcrUjfh/gpR1Zh4K0QrFVDHJJj1lr
9gb13657sVjvDNrFsO0nKk6WLrHG9xqkoD5VOH4EN+mJglMWdCxU4ZVO0YQ9Zytms5PM0wQbqpmM
yI5XU0JGQJ/gniEKz+JlRa0t9/x/Y0/0TCpawnSh2CdfBVwQoI1NVErHRSIq75rr9kSWjbwTavy5
6u7pEhgNb/IT/fM1t/nEfHP60FTT70QHNlCgV0impFs9a2Y2dq7OU28OMtpFiV29L70Knsk3CBg7
XPOj911ZFpjAKHtNjGLdG5gbhzfsBXdA9/fgf0z5xJQ03rRsC+0EENUqCN6zC2xUHrhRheh5qTQE
8KhPQhlLFRDqPBsLA5wciU6FTWdUGUFeJxkgPWRVyEqbBei8mpGNGZSF1kJb0GWFRDNyY3n5CHOX
SbVhF7f2HEwrIXL2d7UpHsFkxX0Cie0z9hKnspYu37wXD5w2tyfloMZ59VQaT6HvmhISJpYIP8sm
z8PGtkRBJE7z2/GXXPRF4rwC/ie0dzBH63HrKO5lyaMaCfwYOAPortSzl0K19oMf/ZUgimKWXDhC
jikjPQmnM1e6nb+0JIU6tjjCN1Gk47oXCAghzNtkJb2hwE43aWuTSnZ+C+i7GFs6Ao70W6dTkWOC
JporxS41z/e0ORiR0vQcx4xmWjZ84lmt020VDbR9bFebTlTAu61Kaqo7dQKr5f1Gnw08NM7ibGFZ
OHHDsGVHaRkT4uQZoqbO8AF4yl0mydcUs0uk3AA1y59S+I5iXeTXvz4qwbCfSm/rdFSILgqIOP43
LLW0kewOXfMuJxed8MTYuQoPjhnGninhAqsIBvbiWGpJd/MwSOJzvzQwoE/TWrjeL15AdUKOv5Sc
vuzEF4/gdLpZEyNg8+NS5ZS966YsgtOeTkdITFtAdvQO4xLo7EtpbyZLWxsBdgyQgMTtFvOHeOgh
UpnmLKlTvvPCjV/XtHCXr02jm3C3NurXmZD39Enz+X9HJNM/wWW7pDFXolqrHehe4whFBTsx0/mt
XA9A8BkjUDJCdzDadPaXerqulQpyH9ahOmFG0S0kQnUUnqfXEm6iiDY2X7sg+idJCWz9C9986VeY
Vxa7ALduH2sMQDoUCBUalzsAAepdKS2bTvj0b/5mE3jM+adqOKDZSKV83w0qSxBE1YBfyJ+A2+i4
7ozuwIq8T7JygCa6V1lzN2fphmmq6KpQ52uER1k+Ct8lwOy3MzMWLRYgOlWw9RmnwKcBaVUBwMJR
5rHkUFDT6/HPdbymxaAqfH7tJ6EqNk7Jsb5LkrOv+aciWmUPaf3lNW/uMFwGx6TFTxAn3vX+a12U
GJmCRoPygcOoMhjBUoxSca50+Dp44CDJcZ3ScAsPH9A1esctjOyPiTmqOyQAB/AAl44efI84aROX
jL9T1u8mwYXhhtvtVhsMjhE4o529yDyTTDueniuK3yOrh1FGfdNtpUwzReGVpibpTojeeI3K60pJ
Qjqq9ghsbuSKpqwur5k5bkPpuNZUPuO7Ss6odZOH4VsCGWDa3vy/T777D/CuMJUkLmeo0rN6KdiX
JoQHNAGHif6nwgf7VSZDkHXoCws4A/b35yv5zOiavFaLlQoMImPjHzsxnmgMHKpV+rBBeV84LIeF
p5PNszy2q7VozuxKHRrMU4T/O/FvPmDQ5nxKUNdVCurewG5f6z73yQygFZd6XBXfjVG7BPMrvUMz
vy07qMP/blJZMMR3qkgMDiMLYopApri8jOJWS9buHlTJdorqg49U4rKbLtcbp+trHasE+I4l4Ock
sRYniFrOMalMnD+L3z9E9WzrB9ELhmEJJZpzom7D4YqMBZYnxv+l28LnWdGHgvSUHGXvfqEUuyeJ
PjnRYKvOWyMHpLklze0ANY9ygWnJDIuPNJRO9AjN2qo5c9+CZdYsdxL/EBct9Yk7ll/LF8wF4V6Y
RGfSTZquCrW2dBQGy/VeqxUKwHwvDWxO5w1IRBVmFsxagb60OtMz2KKDp2hP/9fAtepQP2e2zaFO
xDqhLQOMisWvtjk4v5KPG9Uw+gGhYM72qrUHT5HzVfM6mNeJMf48x9REoKkr4r1oETgK53STmBW3
GeaC9XvdxTp82Pp/f/To8A20oxn/1YOGJ/bBGxhB0nOKIZDlpZvp/NcGCGHHwEXR7oXR6k7GbfdW
y3gDnIlS1u+CK1w2AV3VGrGLGW9r5t0wR/X7JBbtsH6BlbQY3ClNGWB8KxpuU83v+FYeYc7p3Piy
ShM2x/1UrK2AijD9QC2JGoih3DOFDPBRxNocgPZUG/wR1J7XZQoAUd0PEFoSH40Xb83BU8rOKCrE
2ZT3PVQE5NZjvuzWx7XWgphFlFjkq4WNkrA2xH73vnfpaDjRQbRJyLDXVWYIniu3KEQzk80bBdPz
IzeceqxZ+JgtrC4+iv/8tFcj34XhpEixyJOVjjX2pSceroEFqXhlj20hvOPuKncxk749EYG0mFEK
2uRtn0DAaFMpM4ySYQ4PbEYtrR9wKIcDKaFC94QFNlw/I8MlQJrZIkhGt0Ygab3UUtUS8Y25u5Vw
pWXwWWOrI4WOrifh86w2erSHEjgdefPura+BWumLEK50UuEN/PRl7rpj50YTSHgquKtHjV7XFj9X
4V5hDrMcYpZxxmIrCyRTOItm3KNyUEHsNxkYJ4AUS9AlLvPmaJS6zP2odYcdfloM17aQI3UmX8tp
rmr7V9rjzTgdgqapX6FH+chAHyQ25h1xuv43Y0mEIvn/swtXoLYu+3rkHLt7uYn6MOkfCuSDPp4p
aTuknhOa3m97EIXRvvwVMagshpmzJgz9qrtm7CaWuAhnBxdQWPRbppCRyIxflCJOYRadivUgzzRa
aPj5J5UNen5ZUKfLCLgX6TYTT9DGiIW0ZF8xL0V9lKQE6u5tT5v2uEHGvEAMiVboj7SF62sUBXIi
sOvT+rZRitzUBjJYxdGKLCKt/HJ2uAaU1zgRq/DdUwEprpRtP8aNfKvJ0A5wtEodpcQVlUzTdI+h
mrX/jJMnK/4UD44Z4sMdz25+7nBDswAq08Q2qfwhPPpGDpB1zaWIawz5v+GDQx/H4ivFEA3XpUki
NCuqeanaox2aBProIz/OI/amnX1bPd03TSCpgsqYYa+fk8ovgHqolgtap/+Gjn8P9ncr2owpyR/v
Z48liYj2nU5CF8CDQfA8CN2tajnYFr+RGY1QaEgG13wS08oPFcjtQxsIv0buIlol2YR9xRfqptcI
YK8qOmuhw6TCLQZNPGOWzsrFtYJ5BdmMpvIzUODi+TN5CXTVlf/PAYkI+oszzcGYJOy3D0dP8Uuc
tiE/hl5IXU/qQprtragASi7EPNZHhZpJ78MAbR30Z98uIBUK/ppu3W1IGmCTk09xipfXfr1l9+3n
0ylRrjCMCreIR4PYPRETx+fKa8p21dHnEhbz8GDK4y1XbJ/VU9PFSZ8e9ZIEGYXuxgrApNZvZxov
VFvZuh6+OvZxEOFr0WojSZCQE4Dnl/5zPuDTebrv2gFiQFyVUg8uB+1n7akntZT0BmlN2PKJf13Q
yXLtauzTDv4wL0PoVbrcw6SvL5He2qGikwF3/h+cwFLi/itA3vpj540m+jo2MPGbkilLr95HhZxL
k3pxBPG9hZfEAyEHHTHhY3qRbDMuQAGDK+PxdhIoK1rE//iwqw05A9CID1aWnPn6rZezan0jp9m0
lhvoMGjkrL1XfDqgM0zu3YrTUwaBb/IB3TwYZRLqhpDFJP6Swsn4Ki3LbiMtFVwK6H0bWd0o5i0F
VATPClH1SFyEcHDNRaFqha5M1iLM+H7iggHVy9lxviCErfv1g9JZ4nWPXxWVUtfNiYTnVvCC9gDm
F3Cx2yu8hWSDU+QXRs3FhM0piqglPZD2PLfdGDQT29zqIIEpcc+uXzcgB+Gn/To54f+BophuNjBG
Co96SI5VR2iryaa/3KBE5blIm7cGzVaktwZbIDIkTdWiGU5ROrjB4bfXhvxaa+GOlg5hHTaz1ZT1
4UYGZMF01QCfQlGkKmXC/DUBXUHp9hqiikooizd8bpUGPQ2ocJW3awRktwYr9cxLFQ6+abVj2QYR
j8A558xs/Y2/OrzEGrpERRjuSJyxxb8hiuCw1WY0bqSlVeWxdpYuL+8C2fnzKE2xvue4B/DxQvhq
74Y7fv88TD1y0OHGv5J6PC0QGlFE6rB6cr1AyipvKBjIK/K46rFiEJm4yMEA7fbuIt4Yf/uuUMWj
fmipLR89wZVqhkohdBduCt6hDspz+Q2ouTXPYqmiIzlHl+S/cK1gQOUFpwuRIB+/k2OIUsPf+Uva
lRckGA1rNT5ELEBYHrtQA7FM8BwNDdOGbmhWeaTwW3n43yYSgpdVnVc8XPiRWXtn5QxN6+4TeJCw
ETzZs2jzmbyZ7kTSgrVsUODg/MsNGtzskLqm6OnA0SALS/PWjweL0OXkrcvyd7kd98GyCwtEvAA8
gPmOsn1H+FURHol7sAJEkuEFtp20CnNlqwPtuy0/ct6G71mTAC7QyySFiWDshooTh2hLvoOU+QjC
txyOy94Y8yyi37wqVUUvHnlJVY1BmafUN7KLwd/FAG8Ue5YRo6RnV1gVbrYxA6EN0Op/ZrVo5y9d
ska+y672klWoVk9GUhrYfQOHwUsPpm58JcKi9UugEayOvjhjVdUcDvU8+To15ztoUQNPwjSZ6iUZ
pS4JECS9f/KiLfQbXJ7xPS+55vAn+zoPv7HF2hOJMwUOE7gL5pccXM8pjrNgrJNMH2FbN+QzOPVq
Uc1JJKhge63tghk0D3NDjRImFDrH0e/1XSGR0C10xcF93eNzEdDm5KNevOagoNelt/f5eZ/MfS7K
evM2myF5tx4u3KZxBatGpjnR9ngLSsrNSc6jxxxXoyioYxcjSYJqZiQXSPjRMALFOuOukTYTsvyE
iItUhtmccqfPC3R6TQXM2aJzZJUHNLQDDbeqo3apb6O+c8WKx0OhlqBY2tBbXUXMUOm5HzhuHFAF
pRFlpk47o0wSrbwcyRyg4nSQg0QkPSyeQUdR2gUetve1sjg5ScbNYtQAYOU/M8yl8hUBr4awcCfM
IeR34kwnaHiZUabc+8w9az7ZtIiwBAl1XDkxpDqORxj18UaPUY15VTXvEIoWaYpP/KgdWwxXFb9Z
XO3exAK4BaSiUyYZHMbqxtCfL3md75hptYSZk0PCZGSHS/gVXpZ0i/qUd1wurFeJ0dTvt/jCOPFh
io9n7iMPZe2Bl/DH9rG887fWTaiGeuwGmkniLs/G1/ihbiMcHWIfdwMfM15PKSUexuhoHvd0Z6vc
rTj6CXTRJM5tt6dhE43LeJy3A/1QAuIK8leLxeL0OFPdxxZIr/z4dRroWJMWy5A4v0Vb06UiK50E
IFm7hVlxYKLj/793eIj3Eyst5iPp/TusTTzgK7iTcAX2IuQP8yixcQTdw59JMx5iJDjSRLscrIT+
g7kLwC82al8HUHLvYZiKu2DnWi5B7bciMyo1rUhLgDd7LZ99krW9bI16FW5HoTJ0HhezHnR9oYZx
0EJggX6XRBE4ImwEqlAdP+uBg7+RPPgIyt4nE03YAFiW98Eb0RQ+Q4ufBizuxez83W2mlSpmsdPZ
TZ486wItnZ8+3Q6hu4hXWxWor/W8CM8Tr04pJQJUW6ujwyklDBnSzo/YvM8zCk50CyN2aNRBy22f
m6J0ZEI68u5fb7oZt0bTj+TaLI/suTnLtnncBtmFCmIlywM5L3SLjopIK8AvFSMt+5uP4qrpLpfB
DQ7XVewx0i1tVoOTeTw75WsQjvszDdyJC+5NLKQrD/+ri0qlXAyoESpgzxMu6zkYmuFnFu5D0Sen
rdu0vuvR+cUWnux3a6G39IhjygsRRPR1AThs2q4BBQBBnkG3TR796hz1LPtIK0xzJrbGqmr9UmF+
HB4P/Qu+xzG0CWqi0vU6xsd7T89jWeFitWQO84ma3X8GTFYfTb70OfM9GieOzeyos03ZmHKoTRfB
K5xuSGktY5oT05rzYkwv2D5IcYVJ4yqPjBO6sPAhoWy9R+5XhDCNXHW0GUVGmw/tZzQF0Dz4zpoX
fkavNwfla6kBEx04pfK+dd3y6Nts+yhrvl4sX+DdkHILUG1zrdqZamjsfHv/9V82p6a0HHbBinJp
m+IaIy2mnDndX9HcIcOIUL9R/EaKTTxvp57z5fkLhyhqygjx/4U3fALxrkTL0nB06qhQ99uX/kGS
gngxS2wgi65nxtTQXmnDsiAiE4rG4HuWitL87I3E60/jBpmElsefXCmRIDELEE76yoDS4hStzBF5
tiNCnUytfgZ6yPrJTuoq/JB7OyTPxkBDUc7Jb09P6duTmmsWPYQqHBqoVJAv2xjFdehscpLYBFEw
povKi/YXAIIF/W5VSxICgrsYaMUGpwJQReLCr8vkwChO4nLuPsTHUhofV7y+Ix5eNeOgDmPjnuXA
nV317d12Smt3l4YjyngqNMIX6kte7Ld4gcDXFPTemFfk26vBFlBlMKYjFMEBTfTcfwd2OE5eNlsX
dvw3u3Cg93IQbL4E54ypXtjI0enZlMIoviMWqlk1d9cRiwdbA7iI7U81Dzw+80sypK6VwsdpIRM2
Cg9M0Dm+H3swi44cUdSeMjL9ESd5CEjL60XgJMpF3QVvlspJ1GKNoK8bLg4rstVotSNat3/lHbqj
vx4vhJX1+Jjj1Hbw4x/VQ1BiypmBCgW5Jm+KF/J20q/+Dx12YK2wnTC7eR5MPntpdJIsn1poaVfI
ZmCSQ5rqPPYB2G0AXg37mmgsvXi1NQUK7Wl8woaH0uhsGEP9oqqO8vaQzP1Ir72d1Jx3fYgh3lo0
m6dVDl1pegI4FYefOUYvf4yDzIl/+pf3+nqv252XxKoJ2r4hyXDAcogJBArJJYwB1pT9BJ+7pWis
LeOdyiB00I2IStSKzTfwXWJdbT3Y7VX2LIabFTK89H4HYQG32FATFcFerhHPJS3xRT7uPTaaIV1b
t6hj2Pb0i9SX3h8DnnYZ6F9AocPfIWrsPIdvVZuPiXdl+EbbaN+sGrAluaLUEtDljNy5+pMBmzyA
pEZ3EBTWrMnpDTpFxWPVvGoPQh63Ea8KC+ZwLFKTqBXFfz5SZHloXIDz1Bwp6c1pVtZ1uAmFXYoP
9PiAqR4HLAGqRwQcD+r3QZjKdpKFRZzWwfORNQAcWLGg1CA9A1dzPE6/rKQdhBUSUmDOsGQ/CDFR
ZxV9RUs0kIRgodzxKEnc80E6kROK84KNkNnQx0Wz1Uq7cZ1kpD3EiHxSMN2w2reRKC2xqFYJfqdu
hASuGELkDG3QUK1rwrrkZ6QeX+51i/93DkP+t3vK5xdM2ZFxtVBQf6uCfzw2i4xoRSgXMQDFCT6H
Wm7EN3+wkCPLKm7CtRY/98VSE2s2JuUt/LuIOEXWhgYbrhWqhwx9MpqDDBR0B4MknMPSB7V2uYuw
TyTaxanLtuFRFltInjMdIs2umaz1LhJj21oC/9vFTi6XkmwpTv7VT0wDZnadkSds2z86cvziADHL
kE9P70zvqkrBhiYynQxLjXr/jEz4zSI1AyUPjda4xgtgqonj9kG44YAxhAtxoXsL9oaNlD+CANF3
zPeBFYp3ohJRORHKAwmPO8slMyA1s4CVvENL8CJOAbRzDDLaeiFQIVEhFLjgPvwWhaGNduautri0
717vYI3Ve6cr+D2tGP8NxvFcQeCgX+BhOIaGASB+e2v9cxiPnsHY1INs0DNJAxG5U5cISbOCD3Ad
jQgyD8cbzf4YsbHMUmpxGK3yANedAPRSL4RKEgTLVZK+eXx/JitggTiQ2bsrKeP8KuRJi3jiMbbT
3YXiy/5P5HlrbUh1jfcrNgqhrKl6zKDabhyXlWOlASXjPFCi+uGD2xs9Vv6qDK0ga7M9T/vLW+BW
YRSK/B/I/GqQIyzVZRHkDZ5SDPaATTALkRftuwfvhF97cpmLXc7VA4DcbFjxPrVIQ0it4ayy5uzx
7PlHZaRptVX0YrNtA4dNuSalO8lqxG8AFSQoQ62PMT82ojiujIf8TiMMEsiVlwr3BTPcqLknfozW
Oi6eympqwrQxpaULaKTlEI7qFQME1RB1RzZyHqBofma4RLW3kP6fzaXcZkuAoIj1is1zUCd5ktwh
ROafgcu4cmHoUKKN8xVznj+y9jlCspz/weYNI1nIjSGrR2JT50U8mVpgLINE0imIpVab4YLzEiT3
VW63vdM82xWwn7Mw3Qnkq6+e3g6UQQ6OES0awzIZVzOJjWx33vzTrnHHHm2HgC7aPrqOHbKlGAm0
F9CxxjgsMfQG2qX5UmVnVIQAnRpoXmLnlVIRmWinGidBec54kJa9oRDE4TO2ozguXr+5FVE70CsM
99MO09dwr+w2m6O5oCcApUh8loNGTittkaos8iWm/qp1V7d+ORNZ9P+e/jB10WY3T+LcsLQybuvD
FTi0C1lZ0X9MkCLNzQC1F9aw7KpRPGmnWx1+oL/yj8ic5P0dkiIW0Hq6KO4N8wkSuy2sZPOp9ngK
I9sDwDl9lZlrdi3EmtrWEnSOh5bQtU01Scf+sNLsKM6j+PWIeccM260PAhi0znQFK1eIMfbNJ/NX
X9A3+xOxD86WQLRPtv2QSwsUSukJOICfrwaw7DUzM0kHmZKxK0tZVgSm+dahQ+BQkBzcPo/hKrz7
/flxDq19iJSGx7fH/GcIiMm+G0vOVhh9Y/sU2DdGUh/IyOCUmdyMac30bOz4NhlODrpAP/aLm10e
7W0mZswFuR8GkwVAbkm0swGIFj6I/UEI2nPQX3ixoEHU5eLJAqvpkY5WsIeD/O6OyIqVjCaSKveL
zuejbSd8GguixCjhbpbGLnmRoLL0S5NGPLgRXLuB0ZHLmz8pWSoh09ZyDjhUbae1wrIUu1k4eXDP
bUJrTUtAVBFmGxh5KD+C8KCHkR3kmpPTpLP9p2XQlI2N4/FF06WuuKx7zgh83tXI5ttXoThXvQik
lDJqhFB8EtKSJlrtCQFy2WA2s5lZAsRzXGBioiQlFu0dNhSnTHqh/fXQbuJYKRdU6ybyBWDq64dm
7BCJpIwEJypMuazq2mUlfSh+60K43a4oOjsOGs4PTsrJuyWthey9H+MOEYCbnUkSMgE/7fPdUVU8
mJlOublxEcNm9SnThENBnAUxX9Ky2rwS7Lor2KbBo+Zgpc8JkNO7SdL1s5JTV+lFSwCbmDcKbPQN
5suRzWrWvaGMb3JOHzZXsaz6CCxEBeesQTKHvYMZnoVOKuAaW/IPQiydQKT8CXHfKK96IzVaX1Qx
Uyz7k15piLzh0bjmUpU+smJSgg1UnkouGHgVaCNLIQZXN0D4pASxYKbRqfhmOr/e/3szrhOu3nkU
5OATGxv7GPnI/3E/51Gmldt+v5nQ/S0p+eADDhbPNXoU6cIc34g+J0ZCnNZ5nbZzWe7kBL/6XB3a
uMBRNaHINHF9neXzFBavtuaym/CJEzulgIllI6MLEN702gY0dNlYU/bMbhcLWNnZboCf4vxf1xJV
gUlc0GWYmTGMHXjn19gK3mpKqAb5kbVmibF/TftBYvhHrpYnK3U+pY4QaN7bg/fKE+Ay+9rbEL2A
LGItskKzPxrgdRvj5VQRxwR1k1PNGTPGMs9crgpUAxKm2WKNH0jc3mNb96KgDiWWDAw/4Q4wi+hO
jcEbj8RrjTR5ED8GufW/768qa5aEUDgtFZBDnLJwG8Yre0DszORNa0v4DhVyLRSH+R72nqoObkvw
FXj298AGAuCQtX9s8ehwdY1hTcIJet/zyL4VvYyp02iZj/2jJTl9NZiXranunstt+vsr21Y96H58
j0+ITPxjI9k7EA4Kn5VDQ0fY0TodOyS6GkQIN4IRe82rbYZ/ej5ANvhYFYLp1j8hS6h7R02Rngzv
Moq7YIPqbWBjjK0lFy9JjLli5nW0mKDyluoTjNNs0tKQf6N5Aypmm9UC/Xni12Zc371ad83+FdaR
IIrOzQbTC7+jpZ/W2SjPydjEXcAH7cqeYMWR3ht9bHSRN4xh3xvJ5EV7h0JE5rqc++/gScUjQRY3
D5jLdcdJbz8MANLln0CX+9zDjbKPmOYTfINOtmdikmIcILxw1v1HCC/FrlN1I9xta12EgfmqBo3c
twRGXoRVaHG40h+zbBAJpFxXlh+j5ixMZiLs/lrs+cTsN3sElT6fkpDeids/fO2DvrW3zRLdF4hy
HAScdVz00hsDgLWRBkCUAnRHZdpeXDSaKvXxhJI7U1BIaNx7AlBpga+k2CeDBOptFABW9lVWTGlG
ckm4hJprucX8arNjg99wyRVQt5f496dDKQ4IIX5tM8y8AwOjQChxFAFouix+VGMTPxbXKTB1KWEe
P/GIEsCRBte35HhGjEZ7q48zAT6TIYk3IpG/jRVJKgDCuo0G18u6oDvL1I1/pNYdN06wXmbTmBNZ
cdZr6MBUn6EV7Ujv9NOi5zbpJxYbUxcsFPxn2PX/DV31qlrlPtDzMud80CDZHmrxosyujhzsgivq
dzV3+uTSSdT+eD1E1t4kZsMEuY68LkRgGtI6XV5EOGxJhfOvSHYjMJ/NCUVVBWti9BzAUfCl0mr8
kSb8f6WBvRDgXd87zsnU+pGiNVy/VyJABC0eHkkASNJ0sPuzr9TbX7z62sL07/xXBENNkPP465dS
DT430lH9iqNI+xxjPGkpqIg8tb2WRC+CPWjjne+zdgLmZamaCXukqOSZOMTZYdOVXmVe9NZvR9ED
vMiCQM5mbQiy5wJoNtBp8bdOw/jfGXfEp7Hizf9jt4HCDzO4qqtug9333KxTJgrr8i9jT9meKvNU
WmUavgXfZVGo6dd0q5mCu3Jbdss9DirVVx2LgzrkpgufNCxK1LnPkSX+gu+yVtPntup3H49+mGcM
eU/U9I/HljvjRAEcYG91INrg0f/5OFye0ukR99hqVT6Ef4PAEKVwFoFfQETybWzKxz6dBCPl1nOW
Mkr64L3pG+RTVacCcZnUjEXNw6ta+j7p5PO+byn0Bs/ssXd41goRYeMuLAppx7L002zWRphWUe1s
HPjZwKOx5tSYBUWAmKCvoN+IwQ9Z49zopZn99/oq4SvAYglcuaz+BN2lu21fUNHLz6eF69MGR/Li
gj202Ut5sE3nhRxYub3v7jnLXp+/XwV+pP7pxXD1rcS9OQawVdat1IB6pIrVGKaPg1Y8ayz5JJMW
9Dz9/+TGjiMbiSb5LBuJvYQUfaGUkaLlZesbO2adUU7E9toeoUbKg0W7AGsVNJMXmvoSRPHo7MiM
2I/q0oYtrjDqLOU9D2tXH5lee9EvA6K0V1eqw0FCrHOHNRBIXG0h8tgwuccXbgqeNPiM1FcQOPT1
7n1sYWFncSVciw6g07GQyukhH0VdZKpH3ATV1X1YFQuCw3jB/3A9zfAwgTksFbmdY7IDHFSwGdwo
lPlE3sszDFQGYk22rh744copSULrfiKmzcKMSaslcIHgDy2k59YgOF9WsPYdbT857FoBPuR9pkwl
vSTaYPuov9OVYte0WzVyKG80RYwfS35V7/ddUaMsry8p22RUjHVG+EVmGeZFy+Jy0eVLeYuWRX+f
2gPtJF9HyQfPm+NT4GRUfqPpkWwqvqJ6fE5QLlPTrKy0vwrut5eFIoMG521E3Yj+YLmtoKSC6L1L
oWyyCYbn5nzu4YNLMCVqCJAg+OAjLpHCdonQEeC3IPl3jv8yGUrtDijJt5BwuF78NFgbQRCGbiVx
8JrExzmpbhSBikWpMdc5o0Zfvb04KYDCVguDQVtwuZ/HNq5Z3ThF1XXYAiUMrRIBQ1yHdPqPNC4S
0D7huzFUU4+omn3tI6OTANKPZlQxKz4khCHbok0xHA6q48lGRP1OcMIE2CQ8k2CINuVepCjBly/P
zRImPWS0PBIFvr4bOl85tkHkyIQe9Jk9Dc/PGDks/0BIKymKxcoqFHofT7L38BYPxeNi1jewT1IN
DP+eWFlNqny1nvOMhWJloRN5xOFPjiIBvMT4aLzuWo3HYgX4rD408lPUYehHA2NmfJ3pQIHz4FNu
EWvpxG3oOD+EKXINQpN1zatiU26SrLii7grRfPGIcm1uFvHpA36pGhqcEIpAWuYqH8D0H+Vm0V3n
yzJbwBbxlaOGEom/L0PPAF+/fHq9sVL+WEgRhy5ZpyEdixs9+1FjICtfRKXxOXJ6GUKhrbTAwzG9
PVZrxvzSPN5z7fVMsGzotk5eKHk/L9+BiyZI3WgWh6pW6g47Yt6c4rRHlA4elGOrrL5yIn+8V+Q1
Fu7bTJM7O4pbWhSU50TAth3mzpQN+FdxxL8HMSme3qoCo9enj7pxm9YA+WmL+eKgMvkm++VN2XxV
nX3ZvsnU3HjchJK1fRUlVJd6NF8PP+CTcJ3PfnkHP5hKe5JqRgSpywBAxnCVlpMdJKI+wf/hzy7Z
kY7nEFAD3DeYIhrUAXuCosGqkb+rvb4gf6iJ16+L0bnlysksGfX7n/A+Nju1+wJWw9PUekIi1mSv
NGzR1+A3apSFuua0F4m7apUSQr+52OIxoxrd+NwL+axAcQWkq9La2l0kPSRgVOsg0zty+BjZKiOR
FCdtTuF1i5bzwEIRoxuId7b3zEuDNa3pkGGCYIKk0NJjTseCfuoUESOEnjINtVNpQ/ur8AvpAhM4
iwZQjWohv4/Vmt0yINt7MKy1yhMzfQUS0O/AJwG6K9ZUhMzqOVmqqYtANoZRBnYNrQTbV237Soo8
r9ZDil/xK+OOTT8xp/Tm2NRpbnSBExjg5Uv9vgTkVy9o0YcVo6p3WGbVmiO9zfnrAHovASdqcLVl
xUPR4STcV4Zw9LSVVSFtnc1c2i3o+vQ4aImTt92tRBIj5/X7qNr5nm8tF67hWMK2kLWoZmKelUJZ
BFFqIwxluRnTIPaMA7KImfzFdsDuv4wN8Kjq/t/HP5NEGDuFcSDE+YNibcf6lcKaahEdo+9yM+Ph
gqyV3ZuF7PYkMb5Nr9uyy+8WqjmkDKg6WHrONki805QSClO3IAFH5KbhWLr3QslCxOxPGFmT0wK3
CVO+t0cKqlTDg6A0VJVLiVLB+R5SAKDZUgYwzusyhFoYKB4JR/2J4MVR9LOMQk42n5no0IF3nUqo
wJG7atKj50jmEUqOr8gxis4gx1o3AGDHKbY27rHMUDP6hkzJctU3bdpZa0a68gwifwJVjdmN0tsz
5W0EvgMLpWQahFyMv54SNTiRxTo5GseCrIefWTo4X4vf5xiabIMHuaf+qRImM9tW6EKegutSDL2P
kihcYbapRDmvok66X9JkM05sXH2yaNymeuqAWsDeiDoPkf1Jzfkm9gDQ8XGw7OhGpLppDwLuCyUI
4J5l16tQAPUooCUTmW80CiwFJNIofC9T6wbOKIyPQSwd5DdFGR2NNTfB6re5a2xFkA15KplJ62TJ
wmrYG9GCL69lffCpD+ew8SPQtqVnEKBSN57dErrzMMEIFuyzFGZ7Sqfd84o+Lbd3o4MUJdhsMFFn
UU0Jcn9rpzkegxbyDyLVasfs6KUBwUpe4VuYKlH8U6fuI+QPw5xwUFcDDn4frBdouG0ZkSDez99X
N82iMvqGqtkYdlR0GjhzDVV8BIlN1GNPYTxv/Lbkp15Q0dLPyVTYKF1QKUHqPcdLTFZj90xQBv/T
ENP6FbUfxLBIDp0kC7hI1n4PfzYzaNWlaYrBKrMbm+m1YkKRCEzi6nQWehqSwvHXq9lhsFSNYiCa
IaBZ5y9mkphAuQf9Fh7PSKCjaasPgYKi/d+GFYSYsY2e3xK3TlDk6xAkSIa2MT0y5Jmab/sdGEsM
1v1ZTJhxSbgcGZqqphwhl0798lBMqpLkY7N2fMDughb6VVToqjMdSdTNNmf7Cl93n0pLzUTPs411
EeWJS62GCAR6W/lpDATkOrTWXy4JjejoJ+myr1OSB881VjFsFQtBB/OASrSZas7UpZSlHXWR9OYy
dr9XaOpUpr8WBm6QwsBqaxu87VupDYuPKSKkkhRp5U9NXoSR+9GVcsFanQVDn/uYBq3I6M3uW6Oo
s4RCoL1sCOI2gwV83ZQuIf1QTwNTK1zVqdRFbEv8R7HWgtAuSim4oGHU/YcyeBXufFS0GqWBuvOC
EOIg2jUlM5wUhFuKypBjOxwnGpXk1TsOeOMmuSla/H33uhtnjpEKRIoJtagwLFYIHwyjtnddPrt8
NjLAEcj27KNWv4ZLBu2SMK+2nJlUj6qriaSu76vRl2lY3OpdYTpnnBaH+js0EgcrjgDOJ7h5uG6+
7skJdjdCwZnI9/EUevqwiTeP0ooqXeLR+TfsqKh3qTOLPseBC7zVO+fsRTIqcfcrmIHgURbwVMUC
+N962B8f2VcMDWBg9zeTcF7m0UZ6A3SntM0uflIcU9+8Hlh0evJS3yexdpkPmZQOZ48LNE/eXj0z
64/m8dPkvzNQe9k8k/bL7p2p68QAb5bnWhaGKBToy4fO1DLPIvb2PChg0tEgqipA2OVxsx0N49Bi
8F+iO50xblFGcdQQ6ixUwc7vgsQVkcQlsYrbsJlQy/DU6VgE0/5MeSTBho2uqLTVt9w8HlYSawB0
9wj/JgnvQc+WemNx/hQduAncHK+Z+Zc9s4HTd1+61VH7zjoGfS2KWc7Fhe/DgWHQkwhRIt/+AaeE
KHbkl9S4akIkVIu1S6zDWaqSDVu0+qD4KMNl43wB9OAaZVfBSZh3dC432yMohjDST1Fdto/j/TIF
Uio2vEmEJjTVSici8T14qlNMbf59/IeVz3eIu238FVycZqIL8PkhsFU40xMsSR6evxlN4cBdmM9p
TX2TF/LYh1mcbbsOai9WUX78fA0fhjtV4eAoMAQXxaNE/Wxpnb8zQlUHkOcRXD0t0eSCm/HOms1N
tK/fKd7Cac9TvsWctKMgqeINb0cnRm1YvpMIjDG0nHGwHLX20G4ifUR5xw++2OsoqxpUlgr0RBEq
W6klTuHWTG7M57ETMzZ1tA9uv2G7pphAgBQAs5QQo+YJJq6cAMPaclFZti8SXlhPFTjg48O61W4h
mWuGjJR2haDDDaP//vcPqAm4gHeVCv0VlbMJq5KnCCdhB1wnHIMlfXEXjafZxSlp5dSMal/rWQWe
QjO2Zy21WDvgYIkU3RjhAhYoBin6ZlfDqBZ6VFf73hQUk8YlTITP7ygGEFPRCpb33qebR5WmNpnp
0r3cuM6Uz3DF6XOxhwhrzIHcVkY6/YeXHFCwMl+QnuvBj8xKnl1Usr4Bm6gZmS1o7krErloYwZjA
3/MDcq20HGN3fLuyjaf+XUh6mq9ltWsiqZdEiEMCJmisqe0KotP9+vpIDhDViPuM+gKpC4FCL08x
GG066i1zlgbNc4lJ5iF1NQBESrzlrk16imi6MDVV/ZHiJGSJ/SpP5rP0Ki5hXHqaIsNRCx0ecfnU
YkAPTCd3MVKc25f46OKh4p0kn+RSrP6bvk8s9c82yCzpIOdU90EJjBT5hL2+zB+Y9qV5NAWR1Bz5
DRCX57KKD0RfEo6kYLsIkaPASrINw2ISNQLUCpE+R2RvwXGjNoL1Mvz61gEGH+C8d0DI1IlCDqQU
MsEnz9bD8YSZHeReq/uvWFjKeDftq3fM75qPovvYNudexjRCdibkLdZu1ut+TNrf99A/Em6OrE+S
4J/JmsL7WfC2xHxElMQLRrC735OOboRiRfKAsABkMPUD1BFylU11Fy5bkxkRMRPkx648zYgoHqMg
1ze2Hh70w4ORM/jcaeYDdjR1f0qKGhFp1YeZKkbyha4GXrHo9TUyRx8G9P+r4npJ/VpMAL/DTC1h
r/Pc7tjy+SsfvVOKXY7zv7PZ1/JKTr29IOzPsFMdnsBFla3uruWhYKFk2AGBBrveOUfd/DwAg1ZX
FBFThpCk9j20tRia832WhQcy7rFATwSKSrY+pRaafn70nqWcoVIFHe8brxlFQKcKlez4ruOlDuMs
oCfcbkCV8RA0t6vxtdOSGfxF1yt3rorgAVCG1bvDfdYqkT7BLoU6Ft+dw2GjKlIlwUkqXJfZMR+a
i7pv0Jo6UDKujTWog5VTMSV9WEE5FQ0wF2RHpbjzhLTmM9seEUfgRtETbdIfvKrirT9sV/px62qM
TRmneQp0M807v77/vt08KjfwwYEREkybZ1NbbispfIOKVK6tAeID9Iosht5p7ObnRYBDbPFMJ44g
9t42GOtxIdD5FRUL2Brm6PQI6pKODFcJpQZZEspKeCRV9E/XyuLkcGpCg8ntTsPoi8JElCK5HCY6
plXtaxav6T3ZKDEy6PkXYTpZkT0a3ieD51Gvz0k467GqCovv67K7czULVrvKCJYksljzIoDA4pQJ
yPjn6XFy1Rbk96d6eVrXmogU+jlF2mRi7mDyqeo8jOqQpTk0Yyt/XYQLbkiR4crTVIyAPEXuBibu
IiUVf3iqTa8c/z4auVYfvsmBm+MhZlsb1PqHG5j+Mgp/hD+s0qr4lc6oaXPpQ2qWf1Wg4wKqwTvy
9Q6yc70pTD+H3yw4uYR/Ut4zehnxfZZKCCsxuM0dIKZ+CxAIhhqzl6oGB7jF25l538IvjG8r3gWH
sb8ASFZmJyz4oacF5m3z1eToQe1vQ3ZfeBxG/lzi8JAECOhOTsWPW2Dp/QDViO6ftDZYWuh1OFXI
3vJW3Rh9qIcbkM46DnN3OYhs57TpT5UXF5qi+8qV+uoVGGAPN8OQPPi1ZnonauC/sU3d5DSxwUQa
0bjS7xW/NDM4hNLZjDJrP8jfe0GonZITdBhLZtOgxDbl2TLKZbs332QDSqsCAgDG0/KN1I4TA+pu
e5JZ0xgX+NBmaZwcnl7rmpNRqdORM3z4jVr3+VmkeB97VpnqKL/K+2+tT9HYnV0uHQkgB+XBgnjd
dmawTA4Zm36nSxQ+aIO2fZsoqwHnRgHRWfl/8jcbOqki7tqydgRMKMu+mrHv+43IGcFFmEpeW7jf
3AKIlkMR/S0aYpt7wy01VaA/s5Qnye1y0pXmtKnc/CP8G5Lqk4VZHNpYGzn4dXI8+2Le0XQbzWmR
CLl3wgj12uJU4G1XsgQW2NU4VIKDobNOq4bgI6FgC9Wy/wnOqnhP/aiB4iPs3QSiMWsrnFpnTYV3
6Ngf3KuR6Z1xrjyqMWxsn0AFg4iGClCaCWEbQaJy+5HvTtrWbTK/u2N7MqOmmyMW3wlfl/B3IkvS
zJaIpBDUsHhckQvLQBTboYRmv5GxdDD5o/5/sFv6byUjROPIyKoEw8lRczRe0Uu2olC6/JOkxXGy
eLCZ8vKeC1wdhw7mn1XMA0+2YdY8BgDp0/ocQLN254sUEHTpH8NW6ydgp0sUqmbrqt7XuCdN9+Km
ipNTEwOJMHGx4WrXL9fVARQxp2jhOXthi4l40sr9KMBczUyyMBL3Ixisla8U8rLx4/DSKGYXRhr9
dhsCcdkYywgRq1F8RE01POq+apH4laD8OtRtbAsWH/rBTKLTPkt82Jko3qkevm+q/JuQ0j4GqgQD
PcI+WJ4nDQP2zeE/zZdIquCMGAy06np0C/UIo8aslK7E4CCcjcuFWcPg1B6TzMQRohPTm10xjxCj
zlI7hVthVyqXOckv2wkyDXk+nodbIwyxyxW/HMRVv7amEoIfP/n4LJxfWV74p7wMjnRWzCcPUAz3
YKuxq5msazFfNF/46F+78o0X/do/zf9bMp242uSxfDmaOA16kATQnJRGJr0dP0om+Ri78yWYvhW3
GUTSEWbE4B9HYBXgN6ENRLr6ILmPFPcL0veYdRca5hpG2Lrs0cE5CKB/LZH3wogdXBRIgoQn9Vn0
iQjr2b/Dgx+jKhoI1OOaLeeMvBXY4fbwCTeFeY4YYXNuqa2uPIAkWJwraja+XtYvO0NIG3BTlCCZ
+d3bzTvPgCRah938rmMNmw9xqvgM3MOGmmzLuBDE/D8ax3q/a+NEpC4jGMZkSG8DBiMxdra1UDJu
es349dItX0VIamwsZOj00fU6v1nJpzp/gb+eQ9jWfXxG1a2kiTiYb63THb7B5jvK2UOAx31SZ/2U
+wmYQz4JnIHQKAQQ8eUo60qiE2uZhdlBRl0OtoSsEWdQzEEW5xp4IZYAGXDmk+YYIUXen2AnHPyF
Bjw+pzffYNN4rarkOis0HUALUab7Um1v2zY5+FlpnUf1nrkW6u4hVxp0E0ecfzC7VUGHlxClKGq0
aFn9uhCg2D52lE2lSxg+QpHGU3Ae/lMKiqt1gbRW0Ac9m1B67sj1B9q/SkdpanhXI6hB4WmuTsvx
kWNvWiXw0c1tSZ0MUXaPinbpbONomgm+NvWLPTTTue13r/ThooQO3Ba6wzoOAXnJ9NtYBy17f4B3
s56ylu7OGKwtKRVyG1IQnKGgqFz02jHny3uOhCenhwnp9OLTf6IE+F7WllKN5vKllket/4mxVZz7
seGHDh4EavWSgi21M2cjglYy9jHfEE/R4vIZHVQ6zRb7dl4CZiwevjXEI19xhzA0VQamlmkkzkW8
OgujlToISaPQEV5Qazd6Xt9TUIM/dwuzwogEX4SvDrP7OcL11VMb8CYBE+51xUmiAuVnVd5nBl2x
Dg5WrS7pdhHKULnCAkUvl/ZkdvP89jxtzYbWDcYgA9ZrGItjjpoHT0GnrwsE+1WsQFj7JvAsBWNo
+s9aHWyHM3W4aC2g8/JOvF1vgBmtJNSWdkelx4h/poW/fnyH5JciNFHKzopoyIidcVhfnAC2Thp1
Mmo6LgaTFIVSC5TMCoTis4v52iBlxPWORfM9+uVL1ZEzsQnz0VDHVTF3PBLqJbmdriD0eZIBFEgA
0NeYHIba8HQX1CQpiOnUewi3nZqw6WM3KvpH+mjT9FxsCv1SAqf956i+7W7q1PoXtl9jlI8hb8Cs
ac/coYwBaqT7mM7c4/FMULB7keEYP0Y2M1u2ub5RdgUIxHlSNtyISogzXfvyX2ybp6Fv100xQqeb
oLScQt+Se+4Asn4/HZipIx6NV9EfNfNFKwwDlbLkiPeQmDCZfdog8p1HXX0bGb8SOadtywzCcE8t
1CqCUnGWggd/2TLsNwgqqOHxU9K2GHBMo5fICtexr/wPpIWP0PU9BsVlkiwwF/DVjY0VxJWgIMJP
+cKLE3CXRy+2nhwnxSSKDsM/b0kzd+tbGdGYwN02wNYIeRPPyQCNhoNOWB19nlu3l8PUJRa7K0sE
uJ9Bn9HZv1MMHvEYGk33Pn4wWWp4Il4IqNYxn27P75Fc4P12bzXgYbDolrHrZ9DrpxkuhyuMxknr
sr0ceUD4C2gN8avuJN3iivWOz3rYj8bcWUjgXwD8OKV1FmDrOWF22qn0q4f4J9U8yYeu8a1EyvhM
6hSTeGKfJ8+xw7QIens2hbcp/915mJY65/4Zz0Csc3zTuoKuoGvCsbSM+8ik5AMWvNJJWi1e0o7f
27ECXWARoK+u7VHj9ekic7ZE75NqzkPznHwxf3WmVEu49hsh3bmzGSiAjaktT3By2HJRkF8Snyou
JmPbCFf6VQ/x5nHAUYVjwE5akdcHYWU+y7hEkVs30w+n4AiBXA93LZ0kK0swj+8yIWo4HjtwPdCE
6DTTJPK5Rgl4UdYNfWpJUut9YXhvyd8XiQpMhKRDCikzWDsHfBOSjv3fWFlyfglo7F9CIhBoZgxN
tPwHS5pGsgnseZLuwWz7B6+opH7Bf/F2QUBa8CDpRocz0S1knZIMPiEuuo2KV4dRAw6pzP/6mCZX
rMW4v28HaTYwz6zNBgAgwattRQpG8RVX6Cggf8+fqW1Jn4yqDs4eAhA06DTTLheSUGK7hoZtiQMp
1py+WhwZHSUcETMjIgfZMgeDqxFeCwuO016dSWcv4IyDdQjjy4ooS9TwgOBsdEH0AwYzFjzhG6iM
6QOhCQf3tZde3eCjJqnd4+fFmPa4MLtarjtG3m0vg2gzIbEGhxzXshMQL/0GifkbZcSY3VttCUdM
A7LNB/X5w+ZaXbGjzR8VaLfckaNk3mJzYuu3smKkZ8TqbWsfS7Jo6lEM4m9jZWkoTiyFs1nTZjhN
PVjyIxjmAjejPNxWToymAufGjreVnCu5Sq9c2tc6v/of+mwxwNPgvNMkO0rSZD7l9An/CAuwxlvL
hoJPEXBUU8GQrP3Q6RjRAvwc6nt2g62rSSxjyhPz9hwr8Kg2f54JGjdz8EZhoVB8o++5E9bZk43w
qvi8DqHf5ZueBHhOtFJ5+gchNRq1220c9T2ybcVxeZUOvxlDowtWt5mZ+MXaHsbhKsPAr6BE2EXD
+uYCbolT0xDWBYhTRvr+aoI8RWsZgsZe7JJJaPS2EpoFEnqvr4su/s1zhZp1uc5VhrJrgutdjDBm
a6VJbAvPcMhQ+x0KfpSSxmH79jgdviJRNTtsgvHoAl7WBc50VY4JOphyD99D4fwMUUXEh+oRUdU7
nQJUA4YQHHpZZjm9umYAQcDSuS0+CVq3Fp1JD42/dm1J0T6kgzqEg1mOfX5X9X09o9LK/P1vyU93
8NZHSiw7mXsuqnH+olVPqaz2I3pVKtqmXK4Ra8xZnmn/u2ai9awUk/oVqHq5KEjro6qecxXbnt/d
ntjWU3AJAl8y9Cva2UAb2L5O7MVFmHPN7lgQoHkvPGlp+a1laDkhMyDI4z9+nDU5Z9qSwj6DBUiN
eohgEFn/RIJqD7hvVieNr8Twlm+7tdvINHmy5+iw3eEscMwj6ZQ3KldHo7Lhrr3rXAM0+PFEMaTE
8V9OjqLGrynpP9OmkudtOAq7zA/w/mGrHQ99zHjO+z55dWfhRuS/SCBXWQquIHGAS7wG97QXDKrk
dJ+rA7Iw0Yn4qhVa2mnr4FAufugpdHHMqyJYqUYy9cruq7nb6sF47QbXvchawvEffsiot/wMuA5F
gun+pNI0WWySlKK+rnJIIEr8m5px+MXADf/a7LkQ1wDhv35IVGbbXNvb/FQiOgfWJjRvqvBC474p
g6mEiQmGPi8n10JZy7hRIZBAOYcGcNJ05FwzA8jZ/5sJYZCQnYLt1HK0U9mLAGE1BQgaIFoQksGg
ZEvoXiuU77F2f/oMlXW2/bwHqX/jrCN/TMkTZSKnBGYLXFj6sN0sW4t8y7vmbXajfLtGdwtaQJLL
IfMLSAqXtGE609hlrQg+mdnBXVPcoAljj4EjI28v2MJwI3F1wCu4CDFAOFAIvu4j9k2JAptVId5F
4ng3Lyd1pZ3CB5lEQS0fkv+78CwycJXr5kCK/lGyNAQObUyCN72VdNizrUdmZEE+G4HTSnuAXqaY
S0/iMFY2mVth9+6zwpdpnZOv5d9qaFXUIOL5CKQ/z222SylpVoqa52E3VOMF+eX3SrPhtd0HHl+c
yO6z6o31POXMRax+fuPIyEnx8Wu1Kn6PczxGbAsKYquj32esvuk2gKve323dRz+uZHonkYGozZOJ
YcyLz63/Ekd8+EQj2HQDE/lD+6JkvOlRZf2+ihJ+6XV8Bzsf/Ui3I7/eEfQH7UvuXmI4+wnNvll7
xR5A8hWhoRDckPuYUAbtBzIJmFw2KtUVzIfqkG/b9Cmo8HqYNtjLwvL9DnFJPFyA80Km6YUOXFWZ
wQu7uEdg7PTgYKVgg7tEflnzgUg8Z7izIV0z8HMRl0geIs52IIdEwsUjProRD5+jkfiKeTNRuerQ
W++LD/AC/e4tcDdXwCB0b5UAawD3eiqt/OsbvVjODH2iYqIoH9wpeJ4I+oyPQyiUPklxh5YucZ7X
NukJ/ciGAR5s6r4amvXby5px+RMq/bZo/W/YrTqL9IDl1ZDi+LdRBBFMeo1c0ig6CjSQT3ZwCPIm
bMVfiqOLwBHSDuYPNpzzB6FV5MTiZTcgT5GlKUAEy42FSHU9JiUeW+aR5Sea+KKKYMnNhtFpviBR
zlDjIPfcbUsuEt4mXT/nY+qgOZDPN0qN4zjnMyn707eBKwr+g43URQe2fC9o+MDtatLYYSaaDYvv
JxDPo0sTO+pbLLd9CZ8/1xGokvVyM2MARi3PjBMubejgBbhfwBZYNsgQVX+d9iz/WujleOUSKBAp
ZVQwbdcr2FKtT1708MC3j8LnfqbxbruvJu1Oza2jApK2bugczF+3ct1JqNn+o0MW59SNwVOnS7kE
2T8OuAyScC7t5n7050olx2Lars+Dy5RvwDdIjhBeO/rMxWCq5rN3Kvsqk8mpSywo1vEyvjgcnkT4
nuJlE9kbaxBji1ej49/CwR8h9AI8a5q3v7mHZ4KCA10D4Xz0JTnS91LpXOfGjOuuQxfe+O2nsfvo
gH5Lxmk8Uuamh+h7nDionModtaHO76/3Mm4fqbRK1Ut+S/aAtYgjc1r+Ssoao0o4MYIE3b3HqQSs
3EnF3XudyD0KtzzGoaqE0FdSYPeLgx4LD5GF1BsCZlHAZ7htBMS67AIb79L5YuoQiuGK6TApI6WK
EZ4i6z5EwSGEaib52vYWj++nu+WLtDXMvmrvwSLaCZV3VCtWrpJ5SnyQ2FA5Zy6M0Gx23o+NM1PY
fngGqZjk2BrtW+/7RVt7Fneo1lYg4Z6K8tck6iXRcug9xs92jXhSO0w/7/5OrFJZpJNUm+f/Ugky
nDjEO0HTHNeAwHlEwM4wHpt8IVvMDbbFur8qEqPZvMyoRJVuOMNvvayZDH9p9yyIkTm66NKNytQ9
c3HVQOdUiNe69oiXmq6EyfTR8yeqiho9WLsrvhfzemHr7cqbYMcHxhgeb/U9p71MFJMvAbuulrhG
laAroYBo4pv+fESWq2T+7Jbv5DvlMSMxdd8TqJTdyhTaTDGPZDgpLdQXReK8khWaB5tOKwCje1Nj
P/ROqt08yHedmBPhbcTkkzM1LXaLSdj7znXKt9hs6ZAR88IyXl03e2eBX5vbX2zvXkLA8JST4Xs1
edlD0fDzFmdQD2CHmoZNIiCph6NJ6StVVAcbeRxXSA+B04/iKA/eKy1DxBLZiTMiUnffAqMDbKxE
tz1drW6k08MmICZ11PK4o/nuVKrxSbarwxu6v6fPUYhd3U1WyM0yeasgdONPSsTBrAFEi/XYNbku
Xy1TjIzKHIDY2zGGV+30wBeTMoZlKdlfLuiQr71UJCR3I4ERisPhADJVD0hpkPzGz3z9UqILDCs/
7+iXuqfNHwpkr/PXbTJiSM9GG3EDiVr0MeLDKKbB5UtaireRGORu58pIN7w10v36/QhoG0yj67v5
FAv7tMMV2xClKceO7PjHOcvy99PVO4rfMB0EOkA45UJpXBqdpmmwpBb6r4MhEZelTmKNSDanA7mX
qAxsrN6pGNEDxbzfG4AYLRyD6lxYLISCXbWBnIc/B4ixWfLzSOiHoBKRCXvIE/qjkq4K/cblhaTU
gjP/DDeKSIl6VrQKUc9VDM1Eauy5SgNcQu7Se4ZhOWtvJAHw+6+JkKswu3rJDjCoZw14RqeAToa4
5Ac81xg+YU6UYm4M0sFNUDsSPsfNcleQ1N58ZTWSufuYM39Hbl+dkkhByMCFbAtRaDl1y20SNfhZ
hNRDXEx1Q+u95m1qwjxrJN1VuEf3nnLjHqKrwN91ty3dm5eCSaxj8lyMHqPEVLJNQA8gr+njXPoc
oSlVkyqP2IgLbWY2YWF9/t1Lmq4K6KMjUn1S89WTlYfmU4NuyaRYyatiwqb8jLdruP6LpR8uUJzD
HTzRSUzRKuvieAonUUnTU8SQ0YT39yK/ezoEGamgIXW9ZbAO15I+KIALnbm4He6ZGMs97IT2jZ1u
5IGSuynAS6nBChZ6U3wIeZqe7I5SU687Tk47ps7ahKNrhcnhXflGEEHqXeQ+fDcVL9rOf5m6sjIC
mvK2iRMG2KRj2Ry8Nn0accxOTDzLF0SuyXJSzXznw8WTouySP7zVVhIXDXkkqR5VdY5GWHyQ1/FZ
miVVdhzJlqWCbe3X/tnqEs/454hgGE05RfUcPOdGWrKSF8df0B+GSVfuwrIh5P5lFkO9MVz7dHlU
BrkFsrnzFFq6PenmQu45JQdQ9p6Kzwmqm1BORPnOnBMYs4sQHU0GHBquEPnE3FX3Aw/yediARzTi
T106dQRSQgMMyAVw6gRdkAIOPIFYaOv6rDWm++8iMdJfC1K3WganAYTyVE6UkIas6X6o2ssoMWaF
Y1no0ngvwnMr+zlZC935NwvVmhWnPVas2PZPOexWNZaPCGpqY5rOyircPJ6mZykRjLKOkGUUUA0V
wHQQtr0ZlqeCsARRUHes46q8bjHLwdnG1APr4BRHwYVKolMSiqGyBj1mPfw7swZQh8K417auTBiv
o1ZOhxzaIMtqy0Pn+mU3bI8oCnByq9ocyTigdYBtR+iCa2mXe197vl2MqZXgodsjgOOushokOVuw
Fd+7fvVHdv27CoauARITE3wPymeYshg1vqVs4qzTKmqRn31sC0nRLJYNAiQgXBNHpFSlGNxtrCfO
kcdL9y+kAogTikXod3rAByJim0fml6NFd4pVYxG7LYJQIbkNKawXpqcCubZv2ahRtTdKpgdAhbk8
yWtVWKvMpl/xWKCRU7zXsQoSTKj9CXdy0gzWOhpWwVOJD4cWUovXuyVayD0V1Nh2KSYCqmQ0gwTl
ImeBC+qNTEQK/CIYx4AvqWNUZUcUw7pU8ewR9uM62dfqP8/AmCytOc8aczGv4HUkp+UKZUmaLU2C
I5zDZm8W2PWGrnaAJDIi5BNXepNQ1J//s4xaVmlVclhPcR1nEglI8EK4KJ1FhxgLPuTTKvjuhiNE
HAcdG/wMmEgFpQRsi8mCbCyyltR2orr30VSANM9k13kJ1eKGvAedrcTlTW+Pftej9RKRhioREW7I
t4b2ajI0hVxF1ipJ+SUz56qKn9O681nnAuuk9SNAPuTCYnP6n+4pEjHBGejJd5yMOqF3WGn1yV1w
kTH47P6vGey21XzsiBUGzoRhw8bLaK5YjU/An1Bx0L2f8NKpRW5RFOqAoYcnKU8/THEaDF9jhiZX
imjvN+oonwq3Bkxk8bVEwwEfXz47anVAdaSM0mI7BduTF+ektJcogDSLtcs8AqCXULFYJLRdp04K
mGbom2jnKmXK5mh+fryaWSHOG4FsfC/90PqJrHbBbJyaOIsBhIHrpbO8BetGIocboUf94Ee9wsOE
JVLJdfx26bXn3uRDST6Xvm5adfBDG7a7IgJnOr9zPcskLkSVSigQ8Uf4kHfjQYuOwh2S7JV3QNuf
GRUaz+6++KsJrquewkEjrIPbRh/HhLlr0a/Zh4s2I+JA20yipUDmKHjkfmU5BwF3G05/qs0jxcSC
dPZXsV4nutnJAHqUsek4FhcF2JZPEmNz9g9lVKSuxBdnrDP+nOGzozhPNgD550bUVdQYbjIqyhsQ
G26qWQir19UWRsDKFyxt2ND85dtBeWrjBLosWoc0gYteFBvI7nIYP+DGnhW72hyH1iocDQ4BBVCL
n7vHIDgXfg14jqeMCmVomy5VZRP+T4ui9zaALwQGfNVWC3QKm6B6HBKnI1A5EheM6/OMF6BoMP52
879YGMxuzpwFM30zho3V/YSFVmvaUj+gzPTpqmSFtg5jxLxMPj6hqE8whjJAMyLkorv83dbrFncI
2bVCo0QLANzaycJpdnRyJKJ5l477RRL3fZZEqPgGmyuKfxEs2Vx09HeGeddkltWwWWg7MmFKNZ5r
AeSf8f6COyFzOWzRjGP1mktXOth19aJabOvzkhbyqre3Bro1NS5IyXwYQotl73mGZb3OKYj9Pq6z
aPGudrQkY/+JYW5H6+0nCOT34ljcRUiFR8LogfE/iNUqM/Kr+RyiwtswWBKKznbSF1F2uoIHLzAD
0iHwchwz7bOCmvor3KDfar5xZHoO4mzFxlXbOai8ptao/FpxsS3frnQoHKcYvCM+Bflvg8C91c9b
vScMjn0MTxD5Eb5bh4HfOKGbTsMcm8uFXaN6khYuPiUPGuBCkat/79tbL92H/2vFeu0bz3cFHGYg
K3LCfqSoDmvsXvh4X0J1JbvGwzY2y44sQWLhXw551KtotcyC8yJ0LvbMUd6X7jvJ+FyZ/cLv4FV0
VC7EylczTU5dAI+24jKtiqdoLISaxnp4hHrqPkLIHz/4AemMJdufv2QQ4IpfJ7INudMHklXOi7qu
8L8jKVa+PotXYw6LgerzA+kNEJB9E6KkDKyQUDkX8c8Sv0A3e758VHiZs98Z+exM83ki981UFRGv
ikfAB3aEcluM4hNSsOYKg6UfD/Ia3h5nMw4+UNdMmVUyjvJH7mvBWSvpD1ZhtIrv1LYRmaKJJhU9
7BQfvoyeeiEucTreOoK7CcNzpMUPCY1/Ge4sI0cGwhVWy9EhoQZeG4SgTgv7xVEhx0A80RZNANc/
ZKLPq2Bkr0SscX5po0JNCAlqUCr2BQy46TpQbeoXDRrcw8swejjLlWxf+FxlKTa35zq+Y1Q3Klod
wdeM89wWcNIn1kGShBgDRYc2ETr360TNqCHf8XHRwckoiLPeHtbYRxqpyXlgH37aprdb6eEgYgoa
LsLj6uN1NLXJdqCPe7jSNZHpwJJOH2gzu1vXdXUOQkphh8RacgJwc0hPtZ5Q/3IcESVK1DlPusEd
UrN+ZlDtK9UY0pVTijpksgqMBSnquTFFyoiwlmEqllWONsUHkV6NMDS2eaVDO4qFfDobS8BmPf7Q
dUBv/NazeNwJoeBU8eD1pGdoml92ojfMFU4ece2x46Uuxiv3rVmpyP5Js5wJofMf06py9msL3EDn
aFHfuWfHaWwntwt81yS65OHyhvXxVfHmqSuhfBjvo0C49oeM9VfRV3gRcDoaYj97KLQR1HEjdO1I
vIfs9aTTXfxI/mbyDn94FpD93h99OLI36hM6mgoiWsvrubU3whTK+jV5yR8k6/NlCnrC7bYs/3kr
5qpAyE7B2/Oklj2+fIpjtBGgznoHXx4M1yUmAbam9PMVgV8zW0j+aNDm/doucnNijh1rtgoFzZZz
E2MpqOau7dOUZJYQJX0iV8pUvpRl6DEPPyBBReLFaOV4LWhsewE8FgoH7o8LZCG8ogTRShHQGzVc
Ro5LKmZ9XfbCycS11w0cmU78jBXDqo4BMaExOs84uAUPiSWJ++fH8MKbdsOVCRfkVCix4dpy7uCt
LGSCwvr0XMRiiy8ZtEwU+rdCO7LVvO3WOLD8iVqnoOyKYpeXv0j5enPHlM6klEW8cmBZjmaw9KUq
SNGqbMNVlKiNTefhHcv3qrudgacyyhP1thgaLGLdWmgpVu2uTLXV4P2r9+R6Duo5XHuhocZSDg2d
JdXL+1rbQ7GseW98U75yqfLgxC1e7AnB+6CktXBvhWXOCZPK8MPpZxdIUj2iL0i/K1s/EJflya+h
XRUs+sPNjHHz3tyUhaC4uiJPrWDILHjASrtpIkZzSXDCpCS0UzCf4LtPMOd53eNBWylQS1q7tKFB
0yUgsiDSvUCWJkAyWo8LyXkn8pWhSPliTLDcteyzt/WY9qDGbUH8ZcZCpOj2SqcHA40n/6qDtHV7
WUVqSuDB7Upwvd9LQWk7QH2muVRqipt+jQaBleGUD/F0WM8J4hh+o/JRazfr64Eww1r/L1Wc/vmG
iLrgCqWTBsB6lCH41Qyj5f9GdrfKM2ADh0o8MJcWtR6k3rVFSDnrMU5INuzcgpGDIJ78CfPNE0C7
rjrwa2YhO02tKC//OCNXg/NFIzPwTZAkxpI/jo+vkLBlMCAg2+q5KKJ3piOR9yAuKC90NDq4vWTe
7jFjfwnkVZ11Bdd+H8KR3FWT4PHVUGltPdsrGpAFDJAfT4ctKzIXrv4SZCv7ShAW5qkF+bqvvDUc
NyPRGxDj987DSWuOeq8khRXAdPVCprCw+/UgY7mKG3f+Bgz6PizsY/m0u7nf6IAwMzFVJ1xa1RZ8
YcGIVOWd/VZy8OZ5EAMZO4kfnjf8RijCOklpBLmS5sXBx6IKlfj9ppJY7Q5Z9D06Ea2D+SES6VWQ
5TneJlKk5HIGuvRATaJq9GM/NntwsAXT7OHe7jMsgX33iQCwDCndZy47W4af/gUxDxadGDVE3jzm
tC0xsnVcKj9TIk8d8rgfgqE1GdqJELfdmHlodGFF/GULeaAO+vNtoAMojOw+OtpC3E7dfnUtKglt
OTqV3CC8CPVONF6bGWfenNFwSR4xK5mWbrDuFzN2Fds5NkVNLUCQTycx8CGs5Vl5dmM0EG8VITNd
BuaLxpGdEXQSZoMlvVzx4tm08+pFE0n+lCksBhz16EJFiSJUSEjJT+4D2zRQBWZuRQqO0uVqG+3A
Lx00hgJE6vNfZrb0qOyM8EBvidXfSiPCw7PhYZBXYWfWPQsfK/uVdm5Akx1p3xOy6lsYP4qvv+/I
QEM1XcLResPui0PHuLTCdYfPpKWXwdvxasuHCaticLwKOYg9tXQRFFZmldOzfdNJGsMwcxMz17F4
zDbIA5OGFyySojsm3mttD2kaLKKsvCqJQIqrIJIZIkHtzeUx6haBprIlZjseP2DnzA29b2Zly2R6
oSCb2lihgTBLDu9n2IR0BW7/YmaISc4YVS/znZn01B8eYjlX7nCDtOzOMn3NSGKoveYNVAHKC9Zs
Vx7jLI+X8VaCq1tHgvA9hvbvC0TRzopWsInaT4KVcFDB5NfNnbFU+QTCHShDZJzndbl0OROtrGVi
mSiME7lEcHJ0IFOgfGErX52umVDYk9Lu2+93ITA/xz2Lh29s+athZpvF3i+BkTk3OczMkGPEqFZ5
31gAEf/08gA/R54y/7aIKtRfv8jU0xYdCR/0DehfQUd3Yz0/S1JJnTUgb1EMxJtKvmX1lzV+xMc1
7nyaeVHpNZJMSSugS6a0OW9gdFDe6Tctg4JaW49SZSu6yNrOiY9xCB1DYi5VtVK8fS19EYyH2ao7
nSgc7UGCQ1zvxUjo8qikQUrDtpnHlDroRnWayaBpnm3jI0LtkhKEl+jU0OanBMVo+hLKQ1b0KBnk
qGQwCo8c+UB8XIckmPkULkVHc9FbLhoOEz2BZ+1WP3uvT3hVmBmjKh9QrMj2eClNvMb1XzpSXaXV
2FJG4s9dtxYwInt0iI50RQvuU++m6+IBTju8dLNHECSanqaHvmfnOOgd8Xlvh2H5toHsTIojIveM
s8pgQ9JCAq/PLQWQOfa7q/lXMT/uF3u+NFRB6Y7iXgC9Ivw2pOAesLq9U5IAaS27bpvK/BvceTlU
KOn0qp72+SmpTSebZZ8yLYQk6HsFgdjKaYrd/srVNOTo8qAo7wZuNPan60VcYT+G4BVUoCM+CN68
Q/C7SPt1hcIyAcmfBghudf0de9tUlYrYa2QzgZYYp2p8yCkNLZnDYMaeuf36F0xFhKTQeUApknvu
beN9O8Y4s3rLeuGoTPnGlHLk+mIi5Xx32nUWQw+LalcpScPgKi91nJNSxjwzbz77J5m6OYmOnDeD
rjKXbBIjwDivBoam55hcxpk+zGSbb9mdZCnJ4vUinsd4+6MygT7dhC9YJr7LEv1UG+9gfUAGvW3Y
v46t1Ku9klIQ/X+NWRprJZoQKF7HndFW+rS99TFuUzB/42vW9gUrrysCHB+YsQ2Kxe+vUVG0GuYJ
5fEOtZoM+AmTF8WcLBIaLszc/8M6CJUuOnIDXxTN8VuW+78h8nnscjXeeOnfryzJSLVxnUA2y5bU
gqvJQTMgXWeVjCRYDYiESKiQ5R3s8cYzUGL58xtv3DAfu3DXmUSejW0HM1fiWEriPP9pAqwh6XcK
66tn3kZLolL7EY7W+IAay9LXbaq2NMmGwFuGdicG/P/CqDUcCEV5l6jsqsM+FpHvSox6FgAhySNh
ua5cQE/wRooUIt6dK9zJMQYXb0TWr+53eO243lRoVZ77cEyp0sBRcDOkOSkQ0fRXvqz/G8E/da+s
QEPKOt84dpRMlaiHC29Of3SwODoUuaNYaQjRerwO/pT2DKsDlAxyYlnkSEIqTrfCkw58cYGwI5Lt
w32Y+sfZGbdyMRxqytGQ10EE+Xi/2Bunzaywbw1hvE4In1iYU10ywjCKj3MSpqitlljpfejwuxMO
65IGjO1X1aT+rdMfRo5/eeAmiJUdnQ8+ygTGFA5T4SbU6Rlu+UbRO8jbNTKV5M7FC0mKMNCRhenc
y3KqwawhV0o/sxABCWmFF9Cr+KFbUMhUtasFONaXcHR6hY8tUBwutPtCnA6ghiNO6ugFMVmacFvj
gnU2KJJBY24VJoxkctgDu3Pqnja8u9IMCju5xi+xxdM2lVdRRdu6gEYzpD+J/iG9qtvGL8E/Q5WU
HCWipL9scG77IJLIKGNAixMPQCPTt3bIe10XwpvtwrLhs14iRBaQbwatPL2zMrpf1kKaenS3tcAT
r1sZg5IbuD1EYuVh50ZQYOtxJEhhGR6+sZl6lsn/9n8gEuVnGQFF6Goqj5jwCf6ZLfkEvfjZvmZt
7aNBIYYpxanP4UIBxdhKlhPCnsqLnbJ/Xais+/WFvOz0JlQJz/7uqO14I0vCkcfIUVkMdqefxkIg
EtheaDLd13njgQIB409XQVIhoRTywOcF8a4U1FCcUF6W7vH/G6QFeXkIMn/WRX5ARkZ6fFTTqqAV
tQ810EyU/UDVDvr6gFIDy3YZwsGGNbZsCq4dSkGfZ/U2gxw4agQQZ46yp5fC2NlSESrVDgBX43o6
2TWoQghnJk/hIpw8FrD6eujcEMajFUVRW7018rL86ZAjO8j3unlmY4JMDnocwvDob1cNYVX7U9L0
4jTLKb1HcvMIVhCDiWp8I2QZFPDYRWJD5zZbi+8k1tD7MJYM4/LDeY/ikztgEnhzkc65Wfa/EvQK
0bjB7fa+SXnycRTjsjgILM/DL1FAYfhVQ8AJK/6fQiQYmqMdM+CxIfVlhvM8+A+KIX5MdfnpCX5G
lQS+TAGUBeq2amMp1j2Pkmu8mwcBDHXiXJ1odjIhHvsFZNYWBtrZw/mLaHbT9NjS09D6UQ8T7tfw
8JzoTEnbs95jQ/xz5pTOOaT/k/z0wC0oFnx6U0yLZmZYE5YQw9NQtDe4gjMu14dpFAyC3Djl9H7i
NlLEa6svhDPtp17/EgViiE+JXyopoPOLaYhj81HvA1aVzM+jGChe3elxSWHSQoBZEBnFHwPmE9Zz
COrsPuTvHfFnnXS5utNHmwXqmiAbj84GmWRgWZOtDjLskrdwiTtmkIFiWnEJWzMdZnS+axMKibAV
MFx6ez++Eyh0+44VBkvoew+PdijGlWhubNl0CkoMCaxp3mS5S115fToZNIKY2BPkv2BKMIAJQeVe
YiR2gsa6YGSWYYh3wkAW5KyJd7v4N5miI6mPnf2khAI9BlXz9WmGkUwuKj1cFMFg7x0KC397uyKr
Sa0jXy6tkFb/rChGDK13/dX/GV61UfcCpKvc2iwFJC23dHkTQ82khMfPtKgpHe4wPXujihh/5ezt
g+hPX8dEUTnw/gNiq2usg/8m+0GtzYFutqo5NW84fY/xNDoHq16BKCFU8uC3anuTRBHaSZSCQ71x
5MfLnXH5oDNNAbzLGq0BdgL8zSr2fPGsIE9i4gsWCFtHzOXfCCogU8PDj1PikWs1Ilmsi8/9wA0h
DLxyMy6MrRrRsjepQsQ8b66df6Zelt0w6GFuE8oCDdAFuFGV4tvuEzQjFeaahKj7PRkNqYVfJESD
q4LeZEVr7PHTWsmz69Jf5q8jRU4oxCQtz1P9tv9jCcrayVR6Qyfd4om3nVQFyucyJ8j7b4tmxgr4
2a1VmFaTICqmoul6O0YUJlgQqjRz0JLTwacOozFGLEdG0/ISWL8U3kfepllvl+IxQYm+1xfawCnS
7l8Q69hpnTKZbSoBVg4cP/gsIr5m5lAoVRwmxfoPRBK4G8W9ae3JAGG/Kz+uSJO3oFSDWhOiHdVI
+PL3BAuic0QILPnj1b5ZqNwkEnx7PryLQ1TRHSXKie317XGZGJPSwbB+ZRDbkqGwGA4R0x4kEOnj
9W34YH492hxvMJf6PymCaOnhrivpXZZH+voEB0f93T8ZtuD4umM24tmgRA9bM2TUW4Xc+zZ7bF6B
1/uPDrvogBCdc/0mGFEbSRl8+9/6Qgf6Th8TXk3BOo2O6GaunjsgAVO3K5Lz/2WCCVrevqESc3rV
8PWRso/TDfiNUpDcSRMm3xx7h89Q41yYVbPb3ND7Q5PeQpZtz6oR4VeeG0fdghLINORKrxq5Cp/C
hI+pEX4Fak7i/3LRo+uqj0Ms62KcUz1LrLKV+JKR/a9H+6IWTg36M8UuuAd5jVTEzOQEqhurB1AL
kFhEEQY6h9kkZVpDTX6yowYnoorsA/MPzZTyzKon7zEJR1n7IcyT0DEUxozzuBrlxaMEDco+QybR
1B+j9qRX9p4XUjE4xQi9vUD49gvF2Y5aoi8VyGze1756VRrn6e98/Rkbk6t+O1Ex1W1bHveDyY2s
NAv6q33g/JwhJFMtPJzk7B/kEuK4tQwHvGGc5nnTuAyhxj96iO5+5CNHRE9hMFvo6WM+cHt0MFzp
8RaDvbAbkSmIEtH0nF+rb9dJobulsuHpJJCdz/V8dhTrssvZUbGxatqHub0SH75buhc0Or5sVy0p
kbWTX4NqfmRgWLok0zP97kewE6LC1LxLG3UOz8RNYEBqcGHEpLnw3TahUe6s5RAquNREaq3VRHrp
QDuLTtnj61IZALYzZX7d4jI8jY3yDMm5LWJZntyP7hY6/ozsfRdSfsVKP1eVI1kpeZV2K3JcX6Tv
u6dRwbrmjTa4XnGrBu2NWDtmlc974t5Btz0oJ22BjXCsshZXPWPWppvI2fNdx0Z/N7WAKCKRER7f
ubD80AAVVZ5A9h/tBtPE6sH/fSmjJGHOA7BXot5OmOJ1TTNU/gQJl7XehjRprAmv3BjXjHWf1Qgo
s1Bs4fsublLJmSk7Vr6sgG8i9HFVgFUA1wqCuA4sMgKk/Z1s9Vw+pJguxmoClPMQduRY12kvt026
nsONgZvHXi/9jIiB94xa/crg0Zd/RpvpnhvEolup0IXGPQ+Q16WFeZhezs5An3sidYS0/XQz15f5
aGap8NDBC79O2pnBTm12VBXcFqFYWvWY7bC5jEE4ZlN77LobSTOw4bbZiHoi/XNYHzUUJId/TV5U
9lyUyyLYVISQqpkCL5QNLBQcHELoZoGm0yLSRlJWspdSEKEBrY2h5Dj4DBjeZBXqU/EZLJJnUYj3
PLEO7wJ6HqcRbi5u8WL1z5OwTy71e/VItG/8w1PgE2Klic6CzUxzasqp6aSR8aTBC1coNBBJvM4r
DybMi6Zp0vSg7LEGMd1+jAOI1LruFnCAWpxeSSkf7rhppMB5Gh8GYIuXxIvenMpGIXysc/4SPbF7
GrycsZ4sdbO2IxntvKIw5ASI+CkjOz6L1fLdBDTUtsPuFj+Ihq4ptT1cMfVUysGauCnG2pqvr5tX
yqiB30Ttj2eN0p2jSY3Hail7pIpcRetLtmIpLyf0bwzV1Nh4fGVuxa1F62yPYjKa2FvIeS60zFVX
DcGglFBRTjUo/yvpe1KkV++ZQKr8hFWdZGMzm6echnRqpJWi8aUrXDAvV6VM90GffAn69b7wyl8D
PPgNPT2yUHKeXmKhu1yVCmXo1OCagM2J1cP+mJyTmW88aM+VLQvLJvHc78EndSeSJy/HxSVep/x9
v2brcCfTQE8ZYoEJXn5iDM6lWu7I5pypUNphV1gY7u4MWPuVdX1hDOsJ1cQ38Txjt5TxAAlf7CsS
WzEBH7yHywqZximeTal+5JNqjXCvKXIpfb6aedI4UYA6ZcQ4oiUAyISo8t8t9UoOlUbsxlrE9NxJ
pg/lQuDQG6ixTkD1Xwr+mCpesVmUiMFnbh2VWMPnUDppYzXvyOn3Te2EPfvnjAHlg+pJ9/xkgeoE
vX74j32WyH0zVRRI/rsnNIj0OqMRG+BjBvxgSrGTQnC44vTpG4VYXxyJfoWbVgz6OzwFesDBPiRM
WZKs4A9iXY1CY42tHl3IC2rTp7pSvnvIPkOFBSChPcgliB1Nc6KqahBt2Hf7YVG93K10hTRQCH4f
urTXVejbb/hGZA9XOX6jbcYph2JNtSIyTbQgntPdkKkyrX77VWQf3olxWY3yWV4BnxZF4teNTCFs
N1PXk8p4s9zgXEmFloTllMOuqVRwvqzpYl2YDxVjQYHjK9C4XhN3oJS6E7AAFWSQcgOERKiiLjfE
JE0O8Ek9LKwe8rWKP/bVDVg0Rd66waN9EwgS5zdPcRSMd5r0pJWPlzh0OQ79urUDYOp0mknKhzJH
UMCAqfcVUk4FioK+f3HLcYsBgnsI82UQgWIOjzpGNUkpkSR5VezyFbuhsdq0Fm5ffqTPBzx9ZZy/
EKas5OHO7bcPq3ZiRSymR00PADMVDZ+Zjdgf3g/KiHY+g8yNL0fpngyFiMxQvrVSwspEiQS03u0d
O39jHralkXI+1u58mBVRetyGV5/CHtfNr9DUci6xUPft5sDUx1Tu7MjUmWD8Gcel5tjxsW5DFRHq
63QrnLrtPcYP0Ai/efliUTcQ/HnW00a7MT02JYcE8mObUFa5Ooi6huEcE3M1L/x/cRBR7cHRT+sG
u0OEFhV3YlgX5Y+vWnCTxRWbQpiCQkJl/hrdmcfDdcgl3yZTLmDeoaqireZUWgw991zAe1fRbStU
U+FOI41gd57M7ch09svpJ21x2eJ1zcAuLpgWb1YQ/d/FvgOyYwy4L7bTpRUkX0AQPdFOB15iNeVN
RsATWhU15GPbUYfJSgh6PaxoP0DbLuTChFaOJlcBhjwFWy0BiotrRxs7jMGbJ+w6gK1yUryGv3Sn
i21HtSHhFyiYVy27VZoVaSuWeNgcMqD8REyAroZfnvkEQRNMqMl5MYMIrYL14vC4Hyj8V6LtTVP5
3eDNdEfTINsDX47kIq3+KhZu33kgT6s7HIR5TPFiGXAMYTqGFSZMkhzngdPPHutXAQy5Du+kcitB
IIxCpFnnxyTMdraJ61zSZMidWaeokUtJIz0BRZ4CrT/6vo6DQinV13+QTK8dO3r6uAtJNiqhkSV5
lPde1E5Vg5/FYLjr8AzmIA7uRl1xeuup/7Zgt7PDQA4eXRDOVw7i+VUDdsHKhY60bsLpj/v//x4p
9sN4K64HmmpAl3vn/riyCPul3i8Ary5gv0DKpQERXvskpSzdMCho39jZBmt+oldp93zl7Rnh8HWA
4TGVbqxd/P32IZaKa3kpN0sD4IYzDlX09gq8FWmpoLlsqE7NmpK2ojjHF+fPOZnV+EkvhDtAnImF
V5DG84nXU4KPAHsZvtN1WCf5ckmkHK3hUxzh4pG4KV4TkK9E3ah9nVi8dBOwjnblX44sk3wb6jph
IcLd1Yu2pZXbjienjA8iY6AtGyiTgIAlOtMp6/qY5UbD+feHyrTsbZdgzZopHfswckg2c0KNZ216
dAb6DsOIemlILbQUHm2ZwYnq6b3zJRMT6h8jdAe6lHybVRyZdvvljntIXvTvdyKk8ncEYNEje96w
M4cHeTgdVjshJINhJHpxNUdjEtwKVVVFsUAJGTacQdrmipy9Jqhuxkv7fzxxyRuDRD86JQV4BKsh
Sa/EmVQzG2DgavNs6Os0fKkOUDpE+5KUZu/vqv43j0HMcdpz3/peBWOtxs7K9DsRrQ0jCZT2Ru9y
x82kel4ZhGREoVUZCtLjHDw4EqPQISwSr8J+ItB8/Zw0lFwwn2gZ4+XUr0vF5JAzdZlp0bHJ32og
fNgrqvp7fKxuTopEUr90Rnqss3/0vJ+uPHHedlxp3bSOHQSuq3mYLZkMVAQsP+xaUR8P225Wn0n2
48bHYhphxGIJ19qPf4H1Hrw+h9Aa00FGKCQhzGB4E4T8jQjN0ApMUc2VUUI+tCnCCnz14lfDaJh8
33Z/2mVLsn+NUexDAwvm2vNeXR3wPKPySGJQhR3XqVFDjLCuNwBCpUlbCgp/k3LHtT1P8dKdZl3l
3V/U4xhjapJG0n7f3Tn6jQ96qT3lSbld1cbXmB4E6j9vjGhDdR8fNfnMyQiaMjt/8EtHAG/Kb9Ig
PVtT3Cvo42oLb7eyI43X/4qpb/OK1onh8Nop3YRlDvNdkYV7Rmz/BKt+cPClHxiA2T4r9Zc6VyCa
LD6zeO15+NrBSEp9rYNIG8bhI03qienvSUEZIaLuZ4MFl6G/Lcxf4Or6Pmi1bjc/du+8bWLX43bD
9HnQ+K21RTvZyBf+062AcUjFdoacr+3VEZL2pF3tGuPonJjStqe/UYlFDRlUo1K5mZ74KCR9sFeU
r1vkbCUBgJsfLU/qnvIwPJco1EpY9/0XZSgyXjakmpMLZrXMxSBmiJBamwik7NafNvruioKvi59O
YIpxbOPgX2FSMHgwGpbI6Au9EDDra6EWlE5/rpT6WcqrDX9lCwIkBFB2ViTkqXrcCvELjA1u1K6J
87fNfNl6Zfy9iv2967O96jK9NU1gqw+XLt01OAV9nASQ2mU/2YLhjGpEv3Nyeuda8WA9JhiKx+XM
KbFIG+0u3NoR2I+HF8Ih7IyNDBwYonYRJkDB0OWl3C0ZDQTKMhT16HXOnrbGefXzUuViuJ5ibq3d
xcFt8di5h+UD1LRQcvtUXZGVJiOphsF2Vij/CwmcNuLFUPlYYuqjw9Rx1hsdINBKjBVJgFqIDOjK
y1t1QhdN6FjYAw8Bm3DzXpW9vaS7U0xQohkAatdFwpS0BOuIL4tSxW708DpOcJQYRhar8bqJfvjU
qoAQRTdMQE9KWZxfUB2QlkLgQoOXwbmI3O41O5dONQBFXg31a5+0GvQ5yoYfLbdTr4PNkWv52pM1
wMWY/Fr6JwDiecuk09jgdLhrWUxa7sHcal7P66NZ79aWdGPgxpJWfYd2SZDrTJjO8En9fDMHrxks
FYefcANnol3VyZT3IfTg1tnyJY0IKfh0HwrRwjTNy9umMj4UurhOewBx7LmtbvSC6031rkOG+yow
J/iwgSpCXV7iQzWW9gFN92jp/I+ngcG6uyaKi11ne3TOEOLEfQiwQqJ+IvZs9ZLeQIrYeNt6VD5d
f6VMdZRLwQoLxfMGSx9CkXsSmXBpxcwq6m6x35sZLSwLh6SJZ6V9A6XU5X3NFEEo9FYXg9jGYcku
Am0iCLppuYlwWUYz5cAYmIq4O97fnG4QWZPmNptc5RhLp//EKtzLz7KqOipVEoANnX3754yzhvS7
BDoX9o87n7iMgvyvNL3+6npFFdjWwq/2ScWF/vWKZmPO2S0Q0AXdBKr3b7OHnQIxzgf8/C1tKYBA
yFO+52hE/Dv4OVixZAqWya28box2G30uIOopV77Im/cuod26T4kYk/YvuFR1Pd80G7ay/2BxnOIr
pV7y1o2Zdy9PjUoAEUGhIQA5gqjKprdSLAPmCKMZ9D+qN12yF/cVfoJdQ41dVdKZT6vmzixmmOn9
5sB3/a22sPLcC7DDbRfWtK1wNhRnaGlRVDfQ6X7HtZX/UMB7uS1Et/2usjQZF5HDxhjccE1gy7KN
FsFcNbWQWm6CcEMwpgDTsPMZS3EwcNlez8nSJ+Ptc9X4RU0wf9rPkGB5kB1VF5Wuly57W1bs5XMM
Qg6a3quzYfsraMywvn1PXwqHMDXj+4qNUnvh47f+g3lImpZO2F0ZX5fLeYCwe9ABXhXx5419j4u0
SSXdYKujQs1flPtWycrjqKQkf9eGA9dwHhB4qd7TXujrsZWtab3kX7CsWg06qHHdWvdtdJaXdFGP
cgu8fsSb3rNYpL4b9M+zia7IMEUQ/o+6Xsel0pIkG1qDw8SadxIKL8a4RojgQpMPLZ6MeWRy4sVm
2w3NPt9iJzIzvt3IgdDE6giIwkjD3JK/jW4iRQwu7kD+gd8qY3+aNs1u04q+wUfqtIPzth9Y+fO1
k6co07XpcTvcQLJraZ3T4yKfAdUfKufSMto7MjRSNwD41xr6bDFzIl5uAyKtUnpI6wayYlW+KOxF
dk4bGG/qWX0xt4M5RJGxIEOrB78PlEXM2LC9yWDNQRSTrXHSrCSPaY9Ai9rQuAZOt0aBfq+MpuJh
T95+ZoUioIMI27OVobfqMAEsR2NWqGwkUhsKpgzkNVHP4xZH/3McZ3OAnRy/cKPSikihWmxVytgy
DCsJ+7DLMw2yVWYPXpDLAMPl1+wmrZflXsPIRztnyJLZWh0bv/FNr6WWj4Suzf8PEqLKFkfP4HF6
xLqPbAenNxiKdp6TlAYfKQ12fjcUR0mchzhAVEjaygr5vFAtHvrfrG2CCe8D2PcVIU5rJ2Fr21sv
oG4h+feZ8h0ZImrCW9v6IiuQtyD68Cf4hhXwlsHjvjZ+YOa+TOfCwC3lzk8ePx0841p+sYyNsC5C
wvV1MJCjJJW+GSP1+5zFZHVd2GPMmFhg2EeM+m1HhrobMLPjNyGK8sKmHt0JGmmWoSxK34icEI9e
AZlKo8G9kgb8qR82IjAhq8ZkC+QvwbcQdC8xl+RRFEyFssjmtHg0IN7z66pdBbUhf0QEZQVGfi1P
VVC3rS/VOc592SdbcqqnvgbdCanptgCXo+AP/lQnNmXfmQjZqpjEMiWrbiWwwkq5K1oJA58Q6616
KgutOv+PXWEjDWEF8dBHeFKkeb1r11Odp7EG1W5PtS47lq5wq43kg/JbDUwvp4A+jxlYxhXWWTNx
Q3DhmuScX+RwMDJhRAakyqhTcWdGBy9e1/XkbglJIZUOLBID4Ul//tOl00AV1858rC7vJ9n5+eNJ
aOxpEzPgTu/dtnzZOYQeAMzRdBnyu3Qa5yXt6eO+qDx6dtQ0hZrJZilh1VrKMKsJNr6sRBnqlhS2
wmiObtOkHNliq/l0CwEisatE8hbOi/GSBTrvuxOdgjL3WG3DyoFaxZtlQKu9abkNhd0PBPqLvGpc
7g+tQJBONPONGaeZN0+UK4MUQA8lNXwmdBdtY5I4+BjakFIQ9DuSbjhtv4BVPRToZUwe8urG1SI4
fjAP0tDqQNRqx17BEtgwTW9GSP+PyN6VEkbUJ6ug+a+uC/11jSpmBKGXW2/zSPWsoSKHBa9AVg5K
w9swZEvdkGXEgT0Hb/cD/w2j7lWEWZ6wVDfJwnrG2pg/Py7OgYBX3xnKVZ8E0MI1RN+iOw92oqy/
1eOpYH4F+rf9dGbujcXAbvCppinnpNh5boCidvgvlSuu8H55Km+xEiLLZPky1exmpyK0uRbJsZLy
PdYPb7B/4M0E7tOdlaxFXZzyighDYl7R4EeQH/SpBN6n4DoVyesJzDxZpA7pdyMdd6C21ksBqUAa
vl5m+q8FbIdln5z77rucYM6eCPrzwn8c1vBxJxtAm/ugaz1wiheWtZQBDAsAc8Z8Y3K3GM2Xk172
E7FFE9p9EK23v4ImLQnYGoUi2uWhqaMQ+/ygRWwKE7gKcm1cLZLWrdUz7V168GS3U80RCiEeqaF5
qB+z6glKHCRCBms7hUaeq2avCf0gVZ5jyZXLFe0BvgpEA/8Q/FTx/ZjHPXny278cUG2kN86iZjjl
m5dz4VY1ozW7LqFKBB2NfO8/nXG9zMJBbD0myrhO2jfGORe6PPmUBGSMmgNBMJiflYBkTnhHPr0a
KW44W3cnNuJfaPJbspLyxDaX0dZYFTat9MXggFYxaw54Eg6lS9Wm0uK0Zn6dFpWBjQh+rtUake3w
fZZ2yAfqX+ctRP3GueCBeH0IHdc9Vg3elt3osavN5ZMuED64q/fuQioyseVhgZT0e6E7sfPV0HMz
ui2VppxuzDe7C76PHcys6Nyb60UxVtuvFeK0E7q7resYmrefhONr7gH5usm0JvQGf32zW54RYkKn
Om5NoyibKPK3PlpOk0RAQH5btoC4fjdfzL0EHA3Cesf0cOL2pjA082k1SBv5BreDuZvjCXQDZumS
svly3L4R6cjyxGptBopG/W0qLlNwOMIEfE+kZLkubCn7TAzzriQANwE74GSbqGkH69TWDe8ctFXX
vSEuGX5ng5Q8FXkE3PsuAfua/nu4wPIbtTsq7KjE6xijWgarwOXvuVSIEZMSwzGrJgKteDxf3O6q
ocrLsqEHwytfCxxVD/sDrOoBhH5pNJZMbUn6BToxYitvPWLgOF8L2o3DsJ4msFZNUp4BRyUeoEtt
vRPIj8UKitcS8HY2FsHNBATQnxOeheDgPM1QvnIkZQF6y34I0jTdJFRviu5tLqJezus+GyfpQIl/
2YG1mrzxonuuOfx+dvomnX2Cj3Q6vC7iL/zcWVhSAbMeXH2HJFNIBLrBRDFC9deF/Jvas7ZUsWzj
H0r7pdlxIDuQcsW3itj3hdGdbhuglfJ1mMZACjg59J7Q0pB8SVm7IefMLVIYrAfA/dlZ0Bm17Vee
VvrpcQ2he4DP3HEjUIG3Dcg3Usur9U9VJhNvb1eOVkHld7oEertAuEXUn9kXjkhBiExrvhMuTcOt
TyZNEwOvBeC8DTtHTzJoXU62Ed9K6WFI5sHWWcHKx0t1OrXAVmVPdINZiPHcV4WK8/OoKMFRFh6U
uV/y6ax8CTyndxN9qUcGPl1z5/zW7IGXHojSC4EqZtwEAcVqdz/Ym+86wNo0b5rSI9bpRkM4O4HX
LEs7qX2qgwO29szozjLwccOCdxna0osds9hnxg7U/vbzVDpJmjXREZsjul9RshCoqyDesQRSVN8a
eovfZXLCqmQ6csT2jB65AptOYtgg0e9+6m73761pEXzAfTqG4pop2ZnzHSXr6tSDkVwvP8C38I8n
d7jIQJ5Pbyb7w/NmTeaYlFQTAm8fnA5ddIFtWC4Vmj/RawjAc2PjlZRICPOTtY5y97ON2ua5P/wS
vuL8g6mclY+pooAmQmKprKGaNRoARMFYTWqziCPdBUf0tjlqwIoR+s9+PWhM9eVEaqn9KahSN16w
ZqMvuph//b1xYvotmY8oleU4caUsSZuG2rNVQ+5lkiwQS0/aohpJCJMh7bmcUjK6KqVKvnl1Efst
awbOmiiE6dpYzgs6r2AO99+GbehY62qkm/7Upm7r5rZmA4nMIpOBpITHkUFo9rMYmBM8VA4r1Xw2
2GJGOEflphSfQNLRd7AfBWryFJ4pIEjCwYH76x4BwqglnJtSaAST4Ynu/SmmYCZXlq79s8wa4wrg
zxzxuHZchtyLSTQVz6ywJ5hFKhS9FFbySfiyQbd66wDvrY/dHniZ8/alSRX7zHvreM76E/fgtC43
cnZhYil+x9GA4lzVn6ejIZLQYCetD5Y10ILwY14NsI2rBIrMO210aUXV8ZMvs1m2wocy0Cp7mfkG
9T4qabj9s1ms8dPGW9gVTysvy2tw4rvwJm6NyL71mIKvqGvZi+hLbXgkBoGoAYf0yS8+Ug0vbysN
MLc5BJXqzGRGS7EMa6NUYso8GZqaxIBiCJB5Un4VNFoe2T9okoVJUzZjpCOwp3se+rsgNb5Cr0Yo
8qmLimjvp41eiV/2+069sbLEgdjRLt7j2hH05Gf4S8VqE2rcvOrFj1yHS1sK4JglwAnwBGWrAed/
7CUIxe2qTS3jSSk0S4p/0z8AR8clNXUDpntOUalvObwGyffuKd6UbwEXNAO0ivFxesiC205JcrDu
bZbvawPmoMLp4GaktickMzgQ/LS3MsRyzzk5i0rkfHSSD2PHap67qUWU1Jb3Fe8WGsbrEDr4F+B5
nn6v42s9kEyWlo5NO6SygPjBCsKjckPPGTF8zaATomx9aHmnWImEFqGQFJC4jN6+XU0hrglURI7O
hVo0nir/ANjs2LO6W29c56/IVv6rxYWFM6RTmq/BEM21T/i16uIHCuDHkqyeaUgltFrnV7jE5y/n
i0EjRxsg6FA0rrrXnZ6ksMnMG02t6ERnNOCnD/JxPIKt8uBZya0FrmGLnayj7lo2SNxqUumn0PzM
zk+foc5ygYwUy2v2n2gk9Iv7fK5ryO6Qc/Rsh2OgYG86N9m71MDHgaGIyEiw01sdZVjladtt3Xza
79jr7LNzlEeTu2/PbdXs66OffZrBvWYNZHeSAXl1DV5aWg7YlOn1EjdB48o4sfUGIaXjSF8TNkzt
MLJlBJnPzHI/5fwl6+3Cs/HsiSjWyFWqTsBy18EIu6TGqebBr/ywygxvGMGSy7BNGHPwQXEXdfEa
C0t46Uv8f+fF5n6cZAJnI9RnF8J/K2rbDPNGADIXsdGH1t/wbOBf3RE1w6WswW9fkLhOTh/OgMff
sMRzGVQ5v82dJSOjtIKO+LdzrB/WQz412CQ+kv40VwH6eHfJIYjfJlgo0Kp4dlE97v9hnewVIbm2
Y2jh0WBc0czWJZm2bG0PXaEIkKRlktNdYL9KFA+quF0RFyq/WUyDVLSbMjImvDEwlw5n5/ip9P7H
ghu3sjhtsdLa32w/RQW7PsJXjdHVactTOyimq1iuE8/yAg6sOPhJ/DwQuc1x+5txsaEnmXU+lxPE
fM3LKILYyMwqTXIKXCh9F/fc1tisRrpf9oPejS66ZOS8Wj3zGdqq8npPb1JKDgEXPA4OaRZgTPt1
CeI+Le09azZr1Ugebh1gxTdAK0DjVeyoudUxu+jKPYC7RJK5+GXZ2e/iYvFjHtXyOCoAQvgIOXGa
LWqcYHmnwYi+B41mRTRsvcs818Zol40fM1YYLN+8ZmgKOn1H9bdXKn8n8x0k7yZT9TxFrn33/zhi
7xV/ive1PCedKqewBM6UYx4OlqdwzfMJFWpb7OnGv3/TGV38xU+JDnpADXC0KglPdEONWzbX8YHE
ZOVNAqqgplw1Aujk848nPPAnwYMb2t7KVzW36LPHXhALxswXWXr2A5teG08vVHk9m6MPRqe2lo3X
RmWhaX+pavDUenM77PLmCg/HW/IMOWsBHKDQjGecJponiQB/hhQhABQtp/5fq8dVq0ASmDe8OZzQ
nCA4B7Vy4lF5N8Bj42xp5Q+gu5JDtTzunGGtSZm65rFiWyVPar/1GA4m69weSg3r/aYgo8H2yUcE
Ntsk79op6gMFoJDFiT6VmwuV7F/NUD4P4oEtelRz0KlHeLL4ZesViTs31oPWpjfkjUCjTE6Baq5G
EofJVTsEidRscNyD3nRp8wc6gZwKoxYpmFtMuLXk8XVWTvhuQzUwgdaz9u5hMvD4sz5Q0JQuBshy
DWqiFwwcCJxxEhRJjvxhUUnxlwg7+nxdAjXPLFBodS4Y9jOUmTtNozDOwDJmr5gy1d2ugRC0WxUD
uhcuKa/ATDtg5BsJNWjHKgvLIQ+jVZFvvLYCpy1UpbrMkmzeiix5E3WFrw7IIuS1bubxMsLStpVZ
k4A7kJtZpH8aF6Vua9NU2MFlfBiRATN0ZRnkfWDgXrUlHhVjNYbLqOtMi5a8LBGaiK2SQ07Lc0bm
LioYgBFYAtVsco/qjqSgMAKYXS/PmNiYm4pOmzxrFlCOQw7VcFZPRhZuxSS5IqprNyEFgPNnl0V3
4K/7Us6fZLjj7/snKtcnuU3x0UwVFk8aq8Eno0fa2i+VSPPUtF9ngFdkaLD9zBa8HTNXETb1GDXF
/sEWPX9BzikFEOeXYKu1Ec9Ixrq+CwLY6Y3lDUaywxgo2d5sDk5zu7sdP9Npg0iKSB4q7rxzfwAj
glKMxVaMaWJd232NrDxKbHgUpAn9Fahoh6ynGLofzsJuZO8P9E+Mc5ts/l0KhMJ0isDNjZ63vnbi
hoHIIugsYIhwp6vRYSQ5wCVc4RmDOM/8zpMAUpcE5zM1ZsjZpiCEzMab+3kQVOCFyro/zjhkkxI5
qItaaqx9uRhci+vH91wLZJJrkwY8uoxO4bCV51U5mEmCB+9itJuMCt55KjgGd6+Rgz3Y9tvkyHh4
gWWDfL4r/cfJ3ycvlG1VHncPKECoGAgOA62N3eXmAqtjvvt3bd8NVAJvnJ86kbcE8HRXUCnXlsmf
7yHPA/E6dIoLM7M3ZGy96VlCJt4gUYQ5+i4vDjZGEsrhq+ulc/AHQU1uaE5Blk2sTQmcNFhIUeiw
560oKaZIrkc+yx3fvVPLGXoDYKYIjy/tYVzSk7tuCs9b0+0IPEal2h0JdXEFyIrpvSk41zd1TvIT
4RF+t4qTRr71vfKRUoIRWlkBlL7ZaSaY+D5ixZ7XK0dmk9zBD6jSU0+F/3XxgoYOaWxaoelPRfDf
BsGVqE3pEN+dKxH/8S/XzY1javBye+LBnFEHFkQ2395kB4xaX38U1knY8A5JbNEQzfOlvXKEsda9
nIrIdcvp1w5v4uw+5XvnjD0aK6PJGCra9JgVnOjjetpC0NWHGOwIhwtT0exYLuhag5q+0nxnGVRZ
EwE9/RKIFRdG7by4UspI4ZeSOQipNwvrWV0pM7rORoXEtUrd1eYHxBPXoFmz78nprXej35aycYyp
EXxMT47WO1j3anLVyn4HMhqUNf2BBztn/1/i4ILkamDW8Qk10335VIKDvr0ZJJw2V6CS+aGYgVOW
XgUuUelsbGwLa+a9Hfqk6Z5MGuw/dMGqd9NvGACPlX6IbTgoVq0TPD3M6KbQDMyS/KT4RLs0Z27a
IajKoTXdosJGEn2ibuSe/nZ8FM35XNd9cms4DcWCspUsUOfVcgToJapB1QRfsaZA3PcByHUC5KIQ
hbkzhLVvEsWA81KapfQTrbhMkWibKgmtfaT100gVXG0zvdU95/Y/tm6GIaIX/wswDvRbVsVazxR/
FDSkoK7nvrwu0mvNjqcd5uGfPaWdBTH8Th3knULoLrsL9wOt3w6kgIpLihtCeWDYafeh8STlsLIU
nIkjyfzJ8M/Bo3yuR9tfLnGg8DjdpCR9w/0N/X0km8WiYFqDMBKKrb5XYy2bo0S/5DBQ6vpJHvGK
NDWAWevBZAGgOi1+f2LwiO09Z4YvnrbuknHv+L8Y91BH9G8kGbs/mClc/HJiLZu80A2dse5+ZazH
UQSjHbh9p2po7WYrWMDjxRUdIS5oI+BEyoZ8UCmyurIMvO5J5fxHiOrdK4YCGvzppgmcHyvdYhpk
MI1zRuagT8TeZf1hvH9rR4mleJ5l0aqI7HLVKwDxdUZlnQtZQP9d7AhtRYlC/R4aB6krxybg0zby
kDAvGBhMW1yrWBECOWTLfWOU8NDZbOs1ZWC9gp/ggZYC+X7JDIIu5sXcBDWY09RxliY65fLmwAPe
p1e/iWL81JgM64gWCzDfIbgAzNxD2xretcog6MPjhkxuMY5gIcY2LTPCRjiuvSXDhJwwNlh6Gmkb
SnZl2IL/S+N7Q5vgbPale+o7guQbZyyvRp6Zvd84mx8LXKzUdtpRuzXpVopfvem6UxqT0b0R+QSx
XK0i1uZFpRQ0aQdvVa2v5ZOOaemd/yn4IrreTohNvXdTkyAj5Col+JefUCfgDailpuH1yf4uB9R5
c9YGJksoN1t1NDOxU+W2d2qHVczllax40s3sHMH1hLsynydQvGo6d3lBw5/dSX1IPFobZQX2qIyB
LTlPjxjN4plwzbY0dzGpff8uK0Sme5dNWawaR8YuevlvmGZNXPlneeHyx2tHnWWmPyU6VYElsz0t
twRK8QDWBf2adKV+3AqAA1G0UhBdRQJGPymAosMijr/ivbPEC8bSoQclfZ+uX16RTC6HrGRKfKZ9
A2pRZPNd0lTDK+fI0bB3yabMRKKpEo+7hnqTSurYhM5byUAGHcNAOMrIqYKL8WaxhVNMcOFu7zQA
34ilD4kMcNjML1H/TVyDx8uFzBPwnmOpcp0YqAyuedFCFuo/Ai2a8vC2cOebZnvYbVdtsYijxYWX
d8/saDmEub/zBTZg4I/nWGUX/dNpxAUD8xFnsfHEVhR9fWqqCY3YUFWtCdqFG+ZVKsXbgdVycA/v
AWu418GaQHAS1F4qHXLJbRfP0RMPFftQZcuuv3aId65vy/8odRQvY0pM7mPpLOxR+hAMxJU6jPMk
2z4RK1YXJgouCPZH2EHF2g5/gP5nkinUtuKoCA6uH9LBePIXlGKPv4DJRh1UebSqBJOU8ZLak6qh
iZ/42Bm2B4GHuuQ41d8NPA1gbyErtPuhQZoH9OeYOLIhoDBDEYjbQKF0KtPdAxuN1AuinOEKvXKf
8dOIAjrrs6VCx90RaMK2WYTUZ0ZNn3+Hrh4YVq6ivJ5I3/cyUx6pfJ+ngbG+3h3k3e+3K/uIYniI
f38CpCb1GAkDrd1EAfDQxtBIa7phpG+Ki6Av5iI06GcnjxyTyM5jWBqa2NCK6DpNRhUQM7CuBEFx
vxZrn9R/B/jNQzRNe78SG7BbJzUbLyxDHqz3pE25DYWFB13Ml8+9CqIiSLQuBxghhWq7YuQde9e3
HZIxJUIYZGR6mgMaQXKfwRsRF5plbDLuXzvAjPUBpxEP8Xn0VN1ubNxb/ys8Hmb9X1LZQXDUiV3R
ZcYMTzcQOaWzca57Z4HvmOmTYwKAUSfKyGD+1QV1pS/rLqvi8Zgr/77oiQywN/V1at4VydyQ3NhG
j9uL4DmcYDBYcWYaRxtx59LgYdt4qA/mI7xVGPmTH8B8EIz5gFwamgh4dhPzUCAyCVchLHFWiAJV
WnxBRzhsFU6nzPKtc4EWhedlD4xPgTS6Ey11I+QHYtK3cM6BcEDVCz4X1wzQtrrjp3g5N/vqpUQD
1/b7zmbkm4A73xAZ2gnXwLWy8BGSgeqBGI9rAHq4iY/Rfy4S9MafM17Ic9Z7fFPE1TVZfN7ufZ9K
wgJlhEkGHt1A8AgMW9CbY8dt+WBoUqtgQ71bOxXpkQ6C4RWlCsjP5ovqk4wvXxNrBvayQBzG9c9A
aM0UedhCCPAeokDfi3DdCb6TmBBk0hJsarnErTrdbRrygvhlDg6dTy4Yz52i53enrPX2Fol6u8e0
ce197bXXTswvVmbbh24voaec6jCb8EYJBL4iZP06F/tYDlSFJFGTwvqm6dh1pA3fYmbnUu+tFj0b
FsvpkwwiPo3wfuFirF7mM8bmWf4NAbYJX6K9kpf2t+pe0pD9GDt8jG0eEgkSg3TiOmB3M1hvm4Ry
blgeznI/s1lpI5w9yJLbC84KyMvSOvng7DA4Ak8U6dpZ5UO9nSgsnW/088Jjcf3SLCplLA4QDEJn
aLZ8M8hrUm3/hmQbtcwTMeSK4B3RKZLhNKf0mzybS3MXMT0dUKHravppNi+vXf3AvUD/qNQ0SKBg
yTKQJukd+FVCrTNIXnQTaQ8bxNOFT0OFhayDPUdTcMBaK9LhbKaFILqd6lR69K9BDzX+Mja3RtvC
YB8IbNaemZhUoRaDdLZUZrPCrP6IzMRPKSjX1aJrVl+ihbhkgdn6TSQ22/RURHLnmwikNnEFHMJ4
2Fb9z7bAtLw2nZKPY8/WlrroCQtDWleSPqw3l0VhRDs3XE8xOg44E6CvkZxbWFWyZM21zeeiHuy/
JFxDmeiQtvOHUHEQ3VcLufio8mVMmgMnuuAqEJbpQ5iygsEo3Ifh347+vtdhbhyzAD6iu0FOM/Hl
FkY4AzMzjSHzC3VZwShJSLmNW2icLo3PGH9vatBbBVrzNL0CUFyTTVpLq3VfW2Pc0jDNM2TPrpyo
3ihn7aLVNFbwXFZJ1Baxodl+GhDs/DEn9MQDGeH61VpQkfCWaAN8q9W0fsBgV5XbsXtQoyjWt4Iy
I5WHaji2hDqrKkMmipj4O7Znlq59dplAd9O+3airjI1C5YHIGy6/ZBzmFcwC3O2XVZVCUDniTik4
Sb9n9UZJ85dbPZ4oxnk8U+j2Z7Nz2gMecH/Btc5IMmJLNmPQiypDA6fnVg/IS3nrJbluPzIpwwu3
icySllkykkafJ8sFXtFcbcHJcWWIPMc4EUZG7AcNQTzpVUEHPqXOaxWzPxnqEX4Y8DEh0Qs2r9aV
YHBVP6TxYyFKsIxnyTA3IuD8cOAJ6swp+oLBpXsxHHxyYQ9p/RbmssMpsiL3nT5fIkKx37HQ8qnj
xsdBiO9IdMGxJSE0TSrPvWa3JGdj3RqrMXosePGVbvPudEEft6D56MxCs9fmbomgB5xTckzxia9F
5m3QD1KdWaySfHB63lsJXaaey6XNu5EBNtA7mNVrCdU9PZZUYV9CXYwmURj55oNfnPw3drkR4Rin
FEPg41jcn/whCziCyszrFzxzOtQGPz3J5ycIqeA3OCvCnI67gV6EKAjNDdlRc2XR+r6Pjel+sHcL
TZQ7L5x//cTskSAAhWuxELGIRcIyqjtqTw43hGhp74S/17+BZMXhJdGZfH4WgYVhquAVY3Tnxubv
7HYPjZ/RkOBEGHmPQIelma8d+Ilo7LD0tDbW5y9M9kA25OBJWe+Xf/kCce7RCNU5tg8Z/HjKaad2
gtA3N4XokLIzrUpa5dvXHRREbmXM4WX2kJH4PR2NJJzmlIdWL2H2olpqOBZ9mJMX1V3e52mcAb+D
e81Mkk6u/zMdOQTrsZ8Y2bSa79pWGgCbIjsY269A2BuLuTe1F6JcLaLPSUza7eS0EjTKTICh4KPn
nb/WqlUs7V6tkwyqUnDfG+51PNHADf+tFgsH4LKkOVzNQX3p2r0A4MqqnjpTJjJLxitnWFwtLk2k
9VTowB/lkveorrlb2nv9ScnbPeNw535UvCavnuoDnVNCyakONYDch+YOOOQ2nJraf9imPJbVFHGd
1hFPasJRTCaaQgnNW/98cQwIIaToCzUnmW0Y1ZiOuftwaQ/u6eccoW2L8hVEbHfMBQUOBlsc9116
bLPTeRDLwg8s1LqdJemJ7wg0kzYGZiNbyJ73wuKvAL1zSPdsRIH5vi6gF/5Qb+eVsRNZMgS2Ja2i
QjExRSToX/jQd0Y5OVH7kaG62EVYj3RFH/easkQIFyD1wD3RQNXLK3BlLKWyt90NoKi9CBXOEZsL
qe2O/FYVpWLCtcngYwy+LYJcGY5LXvLGur3O+6+54LvDc0baBoS2utMti4Hc9idVJ3b7Vgzvtnlx
BKTyQV2RFCVQ83ul2/JnSdFVRpzLtuZu/cnVKjdzJwRn95oV1mgNTIDWjT2dk1SG55bbZVtDQ7Yp
jUTPspoV1rvvcoPFrS5Dzv7pNucbJnhTuEKc3iBdYwklRxL33hVZSvVc8kBB8+2Ev0Luu639udpN
NlqJ4O6UOLFOq2NXEtAOZMSLvuhT9uIZUNgLgDgVBAtKg1NhTakmVSbX7GxbmBwJ8gNDHov8TKLd
TT/GnbHS7TFO1e2s/yAwj4QICi51X19i9fRiZpBf03ItZMLoODcVBAlR/jFScQk6uFb6Y1dZ+AKa
EggDI5HzS7y3+23Jt06+AiKlEXRsn4Y7YjOayOYPn6WykIzROtMJ9g898B03eyVNzLhMHRGI4LPV
dViSxG8sktIHqjXZGJ8U1AqzjECvmivgsD50wpc1lKnzUlRafnmAKvFJErGwVrTOQe3iZC3wx4XY
K6NNfPJ+eEwhq7VlsfnMv6eU0UFjX3hOXAmcTpth2KfnEATCllajfKC6hOqfz5qCP+YjfsMBivkW
6cP4CYuFbc7C7Osc8P6QPkShhorTYImQDnIRbbBg1TgzTBkJ3W9pDckr6RI1KUppgW8d0dwVzwAv
mkjV6UHXCS0C/QcC4q2n5TIgtMPkMV5OSqrKeoSbfztxxX+0Y5nPCir+Nk/4pg58QInpYiEZjn6B
aENw/iZ5mASGpj6lIyaGObHZy2n/xxZ8G43ustpEYRk/RlnY/pfEdK4UHHK95XNQ5vBu6dMGXQdz
mZc8kGEzlv3TpPfFdM7sKp16+NA7ZXs993g/wj964AZDeV769JLOKnBaKx6lUkZ5tafxobhpEg5Q
R2I9Ag2mmzvRzC2JiVN8i8wF3k4z6VSCb1RSt/6Alv47kxSlQyToJaVR9/dmKwoYFY4In4GlJmEF
bITUFX3j4+l+KquTSuIeWZ8nP69RlCf6VozgmkQ1Emxisaoov5vlf3homFJu/Avim7BxxhbgD7MQ
8Z12uYWnEDNtOXaEHszwyBwAprfmABjImMdESNEDoPo0bTtx8J46OrJgpcbftIwlZl6mrHIDHYtY
lWn8GTzLd8W/+3GPyCdJdA43uQEFdrGI7+rd+CJmBFGezGo/b7EiSu5zRI1ofFBqfgbrj/15EmcM
BaF6/rr+vTn+767fFW0JCeCls3dPh2akkOgMn2JrxfS4Bj5wJr6aRqD2qMno5DyJmZ4S4D4f1YxG
o8UlgSq3Nwki2+fBZ9cXv6yvcQ6OdxkA5/k++pfsxQKV2ZoudRA86rNYsS8nzogTdCb8irolZ9C0
5e+XMVLQ115tNvryNo/XiXV2qKjk4UVYgZrOhx+AYZnpkhT+uoVOoWQu+9E00Txs/gOhG+CJGqh0
qZ2mAyTAIx3w4SN+587eJdpa2Vj7geUX29mnc3BSWTxw5TOIZiyQPA69m/tVQKpPSqy6R8WKJdcI
hpiZrvNHLeOikyrRiiL3AEWA4V5yAP3OqCIWd5Ib4iwOsHeWVZPIq/xKdFInocqPNlT71QZdoZ9b
5gCwOFUb0Me9FG+Ou8/8iAErO7kSPPwW3pgpzEPeVLKjCD4kCD3lh8HkHjBdvTiLI/Tb1g9puRwa
PJRBf/S+7fbK1PjW/uFnoVn20Sh6DVgbzlq4Xb6QgS6xcNyZCICyfAn2LvyTbKH+v5qWZokvdCjR
VbvD+x0oMY5i+r8+g4Nd3AF735wCqkhgof/M1ygDIJu4Eo9DbKkANn4H9CQYx7lr/EFDd2xWCYBg
94rB2KgjMQrDFwe/0r2MLRPWu/i0g1/TujHpprb0/CJ8vWDsjt7UuTLVSfwKsxiR9N/1RNlOJHZa
NhyvRtS4JEZgn+o2lJCpuhmNHjYkh6D2myVD/WrZuBUeFVMyjFVx9EHzG44+nAZZYi+eANV10+Xw
qB2MPd4kH76AUjfSdUuz1E1V3U8OfWrDg1VYkjQSZTfA0rEccp+Dda6vAt2oN+QOmcr5xUM/PKSc
oV+s3JAXY3UwSLgQ7fFCSmHsagTaFfkUeMfRMR8zvcu0fmgC70gyoVcnpvlSKH8+mJXwg4uakFCV
jNbKxr61B3HnRK0IeCWmKr70DgJIg7bBQLQzkdhrsg/a2c9wGXsl7D2s/s8DcpqPG1ONOvd0w2TW
6YEf7WO/0obp0zqGdWbw5tqnFBsGubW49a60/fBLIVxqO8VgFy0COzS/zBIvyrRpuLnow/p1nM0M
RTk7XZ2QF50A4/HJ84b6V6xYsEuwJQQNyjFrwZOg9KqTpiR7+tfCSqdgbIeM0taVF+f4Ih7ISLHo
SWXoujeYDzsfiv77RlMU4SER+f18XMKCHM5Wz6RIRcVsdDe9c4793/n/V3ZXSDkhbyXFzg46acyp
aFhjHeqwp0ALmCcFOYzNr+iFz08o0wT3933GYxUxTN4ohfv+eM3PG+fG0JUAS8tphNvyFfiMkTib
hR8lH1vEURTS+zygopuRZyBblQ08qsraVbsfUubY4uSev5ZwgcSWh7YQpV+eLO66eogdIp6a7Lih
4aUMWEUw+eFOgq5n2q+REeGIyLcQ3RHXkAsZKOFLhffwFAzK4MD8ILXMK0GQjArnbLqVDYTJSeyu
BuqlRDYUmQ0AIH17RVBVO0bJx8oghsXuGrcD/WBQ0ocgIpB9McGexBVkYA/IyO1w7MkmMbrXLE3J
vdqStpULgSfzzRdL5AL68HEqz1Jy149IzK+yHq2byaBrAxNe+dnokYL6fw5hLNMo8cLGRLgXeTQg
jPj1Sbaj4zNqbjwRZf4KaMMVc1yCWVe8OxqkQuYptrKr6H3u3Kcajd1QGjCz8GCIW1ZqUEPUbOJz
X/Nke51MV8Ybnyt0eFugQ7yGwB7ztg9VWecCMf2/4KFLe4YzjMVOTUajCVPd65KBzpNj6j9mzVHP
bZQQoNfXNWH7jP63YIU10z4/SgwCzzSHXn/4IUFv+6XVShyOqZWMOMuxPMqpzdxfbKyq1MTA1gVo
Um76cWKOl+v2EcB2SImr07Ord6PgeznMe1F3siY3zuwoUabe+NZ4yg9p3vnS60dXMNRT6ftfzH0Y
8jXajDO1iQjT4v0wf3oRz0zQGZG4yTyl4iKwntAN3AthH86baHMcomUNt/VDjkstBc1lvXXsC9LV
2bvnr87IZhK3HYeZnD6zIZABk+QTWuQ6e1+GHX4naQdShcQJC7SfgdigRx6kx2vrCgoX9M2qn9Mo
iCPsP9GGOyURlog5qUU372HwzDElay5IZnWQACk+FwwSkPAkSUAPu+g1DOHt6LME4+3aqmwZXI3E
zpv6N/rM7Vi/KK73NSeJzygsh1T+DkjOtWx1TJOYZv4IxDjHHPEAkrmCMqYtaYPQho0x+Rx4kYAn
6/XXzo/nE9zhpJdaE8/u5ra4e7QGd7gqAGmrMJqZQ77ZonGxpq7i2f7OrfK1FomaStccLvATEIJf
klVnmVCs6k1Le8lcEyZri6paDPm4V6eATZyt+LbohQqwDx31abzueCHsqyXo14vooisjoY1LcRKJ
XJ63aPyRdjeil5+vLPhhBbPiyMf4CRhb9giXXkKME22hEY23IekOITJGnGjUJnBIyLv6IymMfe4F
Tl3bbpyZ5bhmO6zAhWRvX0ej1SLfPvpqMfa834qmGL8ZTbUDJbAFyUzGdk8FqV0JR16G6xCywcqm
RhT5M/AeguVUf2xvY0FTwgrZwSnb2lYlw730KnoWrfHEk1MXhpMGDhfpLrZ6p+JrDGffzhu397zx
pqexMXw+CyTdv3VZbkOgnRY+VcT53lPv/ctorl/m34ZEofwHCpNtLJXAKtvmJqi/cpWv97rvLRfZ
6rIxSHz8Tpgmxucz/3OurLjRz7VNsX0cLTQmuQLAFO20vzrrmygJNcn40ADGslLeNuxLzlE9JH5S
k2l5oM2lu/TFUKONbCuPdX4d7ay861dTJWqS/g/9EIrPvF9d6V6hPahaILcqNp5o2Ksy8FJ+Ija3
KyhctDrXSZfF/9kkfkKQMZC+QYy880940iLZrd7fIMcPrOMvuXMwuAYx7fNCzaC02VOOSeNr502e
MriUn0iCzxOtJWV6RuGDM1Hv2W/Y8CP7RbYCMSISY55y/+8BELjeRCtMwuy4qYYZOsnrMMl0PPu9
gZZSH48TZmKK2NEiUC2JaZagKhVZPbpjbvJ2k1AAtlvn33/nbznvFyLTK3EovmfE1kiyTr1Sdzvw
ZunhF3nTyM4BCkAE2vYSK5wjUKo9uHaHYy/7+O9EzRVP6YeUeY+QQk4ahSWFoDRdpZzy7QtrrjPk
abV7n7Lrv4PxDtw+m0SvZdPr/QDmDpllRLuKk+hsU7e/MuDJ2RoPQtgHiFrUVUmvnoOOgP6hW10H
gGuO4rInuCvIrWU9b5dNKWF+9Pf4azDxw3ZM9FVx5dvRw8DWhxqYfccLqyBnQv8QJAufrKneaY5S
18dbAJ0OQVuwIu6LKtgPhwOU4VFThZplUc1LHjRdwb3YIzLUuQzWyppANqcEVp6E3D1NUv6Vf9tg
T3r/htgNINa0UUMDdTdrYpGBZibdB/B51MVz+1SqR6gap5tkKIlYzOwJk6EJaH2tVCXzi1Dgdwdp
PK6FWPkCjDlNbxp59WVD3V3AxO2ZcCBUHcrbz9uAg+NTS3ulc5rZfyBUvhkUPSyFYau62eVuv6rF
xwmGjkTmveo4Vup8uRcFP2PQH9eCTLnJzy8PhyaVR0YYKUNTn0I+32CP8ZVgFktKHBT/L2EA5dpj
y+OVOKhxzfE045Fp1RU0RLbxY6k09QpeES5Dsu0aKEHXnbtUoDJbsZmJO+ihoLx6xsefI5Arwzgu
Ta+iUVqd5qOEZaGBwTdMyu2XSfjvBwOW36gHzcngDq/juuCJ+DvbrfwrCe6BCdZcsr1ZC8PvPTeX
3pM4eNEd/VUmLObhWRcCcZ3KwOQLTULrd99mnR3s5H31ZtM7+LdZTBt7BvhKJjzI2DbnVlxiwyc7
EHyVnI7ACfUru4Gf3wa06tr8rSt/2zyPO2EeZArPqenrwGr89nGPvwUhUJ1kgWIzcl4FXOyUsham
r0b+qKKe2Mo3qYKTZ0AB0vnBYVwi76+yYiGV8lXn6hRkZvfBUV/zagOU9IpdcbBFShu4Om/Fv56g
Mgzk9aivdnjYTThH9Hh1DvUm3ele77P9RulvHJvyonZEg14AP6GFwD9pws3PRsohBe4b9zHww69x
2g/fnW8/bpx60Sp3lf4uA7xoLN9eTtK0lrsS/XbJX5ooYlOmamRvXw9ZjQPZ/VATUEfoGRdSHOSC
4EpON/Mzi7p+kJL2TIUoHJp7IwjidQTf+So7JJb0RqHSPnSEEInFtBdPX+h8GR5JS3IASdrvrcU2
F2/kY8y2lOnPJ6nT/2+2CQJxYaBTIa//GGFYT3qrUQa3sHcGfU5gDxIYjWHMUBXP0rhjbTXlRdVR
AkdxdbPlfF2piT7VtqoHYj8NzqhAKYIJywznYKCsYdC2VHuMZr1kVmvRbFAOze+G7zA9PulM2VgJ
oyHkFMCuSHOZpFCHtshp6XeYL5d3FphRxEBTshY4Cg3qHMSLX5BWMfBieB1epd60pSS3nPxOXpNQ
0jq8D0An5yCJ23aiE4VjjXQD8H9WjCslCoXjWw3W8gDpFXmFnkvsY2tnOGQ1HQqiuDyftX9G8Adp
l29HZUZzWTzIFzt3vig+p9hmYFS9ytlA01J4TmW7zIJZLri7q/4JPYHlXYj8dmskc/BSyBIxJGCj
+E71gv74Xzaq3tAIz2yZ7u2gkfhDUPPJVZqNUehg3GUWR+MM2GFsfRfS2ZSKzbBPAHXlWHrgauSM
rNKeI0odKu//iNEF/RFsw95NaeIIh+LrJmP6tlKCSXRNeSg0+IOcd7nlPY9cZ8sQuHOqJWrEAsf5
eOmXaGsjSYzd6Vd6PcmT0Vb0Do+aGwvH9DSTKuaIKSGgKOAasAm2hquLaq0k+FTycCBA6e5aJQse
QFPwzSbqH12egAB05Ki+1kAvjR/7GoY6AfEN4KimxgroJMGDEoutty+b8jGMisPVzpUdHbv3Ngj2
pkwptTQMHKar3fGjHAvFlg4H9q6f+pfozfvNRgyW4lix9Q0Yu/VYt70DIGC+A65T+rXSWPZEecn9
AW19nNvyQIoDSV8XLXBySIz0eyv7+UELJodPb8l8FV49YwVX/Ded77VIIP1Eu36LwLOIvhSAWg0l
6qnHPZWHR8xmOcZQKeIneij9QFApBngblWYUhwa+GFmkICjK/Xo40pscUraLwRaZwI6DygOLBG2F
hTRFr51t5CCCYnY+vbwc3S4qjzSZyqm28NA2cy4jRpf6eLlgzUEwIw3mMOsdJeEYUalkJomE/LbE
S8W4Lnwlwp8a9gI65RhYwRV5rpCEVYGQrj+WdD24kPSIWz1ZBlp0vtxlE9Yj7ygEFQjsd3YYjdgg
KmHR+aWR0gCeEPbUcp3jDms93XiL/i7wdaEwFlwS0gJ1NezidwYnzKtY95zkI6Rnxb6qwQ+k7xyw
utJ1bVTOg+tljgStdI4H4azZy5lquLk0NH2iP+5Qy9IhAQ7c5YoNahyrJoW8RxbmNSLEOM3jxshz
lJ7/SQK/w+V2sKyDpaDd7CPdIamUfvHJL3CupXUea1eN6rXJ8d260fneFhraLH/8vfeM4JZTPM0X
g5I54mHkzQn8D7UqUz8/HAcbqmHjfC5qrjnT0Qtaka8ZIMqOR/ImT7AqNNHRKsA7tNZMLUEAWwsB
pe8t/mrqIlwDJyfcJhZTJ9B04P+zWc2iJqEqAs3Hh/IQN6jo2fBHb33VnJQMSwyn4ZDZ/LKxRzcX
sRj5vF0pPBg9XZSSTeUFeGrvNlBcnRxjvacpeXaLEhsxPUKFMpB7mGcALipG9yHQ/JQin8hJ2dNJ
OJcHxlHNfnG/cOB0Q1fGRLRYC5geiDl3GZ2zMHSniAO34BGCUQh+X8DhGjm3Ntzf+2wSl4OUpIZI
jcs+RXVwz6ecdEkxmDwtLKCcE0fxPDB2AhhAsE7uub/aUyhHMLaZ2oEmKmZX76QnS2uCh2vd5xuC
fPshj89fYZYGq+WbvDYI4GOy0H+XJ3Fqss2kE/JA8CYjGRKMB45pDAd91rXr4p2GP3wwjj8+PVE7
BBOQvhtigrkuFzPodUkhPa6IyMkhi0kv0nDsV75oxNkESnJHJIacrz5+3fs5K9eRY2AwcnVTgu1u
2bVckTLyN9dALc8AK+PfyERHZh/MZMNcGgsO6wMJpNcUNVLmAoCseTjK//pQ7ZYLsVdIOGbisYTB
Ro6rpNW0Q+a+hREudHDIBHTBLQapW+Rr6hZvLrJa52G8TUHjSv6AI18r/+FYfM9s1x1kFdPOcrvN
jO40khLlpm70HzxhQsyMB8N6aa1rVDR6QR4UoBdqJKYdLDYaeTsKK+pAcfrpe1GvBVD7WzLC0vuu
llCTCKzyA7KIFdzPpAGWbTE5dMhhLzfUFxbZHo1y31VqYi2IsDuticcbvevX57KYP2yzkD7MfJQJ
f0j1meSbm8yumvB2qtdc2qWLsKO997Dgx5cJIsQ2Y0AB5C0/hMdf5xR6XtENUU1JgJMSv7Qd1qTg
QfQ4+98MR6FQurj1P3A+da7AUyKlRcH77WnCaiEfnCJkXhLTx1LCcRPQHmdW5NaY88pwNzYTAOIx
I8dP6CE/vYmw5Ezq2NiO4JuU3vngII4ghFokaVyhzNvbmrG6UV0KuwcZi+BRaGRrM9Twj2YdvDi6
Y9CvQS34mqniu20QpW5/GqpT7BCjyp39P26VdkImVzx7VsFId2wq1OtCd/faXUdaplx52y6UY10z
a1VRRZQvQ9j0i1zmVrDvMmc1w7qtl454kXJvkir/lr8LZqf6facipaCLRD8g0gdeFXKt0ndvAsni
9wsHRyAE8kxfJ45hpY4LSBQjIO+U2NOy9Rj8fDwsV5TmGcWdIOT3YToKc/RDyoh8XSG9QHfLZk+S
VuTj1e4UafTyDuTrMOVGPLj/p04xoQiq9dYKBj+uA62yGkkmUy5h+eLTwF2iB9beDvgbjBC0ItP4
5VuvtdArgHIOf4bskrcU9ufBKZXUneYhpnyWttrT0+1gH0OR0lY1TKnG304SG9SuVZMBXrojdhAb
NTwLhZFlx4fqNk3vKQ+FQnWHHNDDyTB6lowW4eQpPflJlEZU5FVb/Icie6pe7LGZ5L5o3EBh402a
XVrstyyjZ+mxbH5kOkGlF1CfvDaFY+7T7u3afBATa82TJIWluWuhbqCRwSGgb+P1am7Dznl8kfD5
5Dr2b06YmClJgzd3wAd5EqZTvM1bWq+X/4DUGNm0+jBM1efDBGs8fitFoF8SXNLfn7J+E7OuLNxx
UpNPbQdw1FIGkCTTf7lWHSy/xHojdoIwAXwfjCEcv9PmxxqBs4JpVN7q6B9/CfEwINF9brYZ+tf4
kAU9N/t/UdXlqXRfqrGlve/1GoJiMKgKfAC520hGLF91otln4XFXjcva+daBcn3vY6dpU7s+ETa1
s+fKXVt0nHN3kUyrYBGi1alJBZoyEIg/QVqTDh8UbXrbv3dICC5pfjMFl+ty0Gl4orA/T+msYLci
tWmFnY2d9JhZjbYL5jbgSvk6zmvzQqWip4ibZ5sU0KEzm5yrtFsa1GC57jQsn/YPPQ2MFXDfH0/s
OcaGzhe9lVJox5G8NzQPimcbDw/YxKJS+QLulIGnKbdxQ/xNi+wYktMA7oG0D9C1WmnwgI+wmE7C
fQxNubhf3dk8c/joGLgNCQwrefHqEb4hNvFqZOp1uTTpZ3f/W3wwcWPqPCxCXUdZXpmNZE8D1MAJ
BN/wPEni0ct0A4Hlzt20jQo0NCqasf1fZVRJ1vyi7Y44Ux1in/TJSpICy111FDIganplfXXuY3V9
gq2p7gq3Nu4OS6m3x6C4vj55LAyhhY6N8zqANw/wzC0X4jf3t8XZj0q6kLxFdBV886x1I4bur/cF
gqvXfm6R+efZNH9ErRE//Q3MBoLMPwByOjYPz7UJZFI79T6arcJLwzx85/EihShPc0P+o99XYfSr
gCmWvHD1URh1rWcx6YHQDg6JaeLSkuN4qB0SQhQqWAPlI1f3djJv8OwocjUVY2zhmltJynujxRby
ioZH8DT3q5hSYruVpjaRuI5ySqhs/iqHSRMTNGdIoRWdTMIeL3Uvobt1FJp23hPwEdCkVgMiMNwT
lR4KFg44DsPeqbDq3XWMrUEk91V5Mqfzb0mnR97m9DvcCrY8NCMSiNQlh8QZYe7dqckq1D0RYzSv
ERr3caGXIhk+3UJd12CyTKWvNhA77bpMk/FNttB8NxtOdy8L9xh3KDiPpMkzDsgXkm6Nc8CAXJNA
AdHDb+YV3aZwFmCgEpLmkmPO/y9Eyg5NfytII2lnFDrnrxkujrGSEXnDzzwua+c/ubfKDUyfBd4I
VnEda01DMbR3thAV8+hZOVYYYZKmOHGXmwMvR2qvhJh+tdBUyT1L8M0/qgxFaY3lMB5Zzr4kVeii
NYs3N+msucRu0TNT+7fYPrWzYvlkBcvap8RIbnjhMkEt13khPTIM4iqIjgb313Hld2JXrF4QIRP5
VrAx8oD9F0ruuOWbL90QwhJt7sLJad9IInqBl5UF8Quop03fKzW6U+n/8tklMN0/0TaF2DiyHmWa
fjgm81Ji4yonGPYql80Vz9v3krB+H6UY4Tn6UlWC4ATWU7byHxBbYExl7r4NwpUIDN1GeCe1lSOK
+aY4xpBxT5A6vXGKfl3tJBzpt/Qvtin9w8pi4f7i0J2Y2cURTS19kRVkrB5rXqeMDzVY9kh6d7Vs
SugbNpHjLU5GggiP3dBRj4DoS9QdDndsHfeL40yY7kuNt5YGSOv4etZIfQ+NG2h/cKLyM0Lahi+R
ljDmppo86p2VHmEvCbctqx6lXRiJaOpg+6Osa7VVp8uuG99Wae4DfEwDzcuOtmyUvpr4GAPc6v/B
BqsoLHrBDVdlOv99lX33W1LVHdCP8flBL4sq3RwoFaVMlw22YDsu3t/fvolQM25qRvzEZaEfZMQq
2936PeoR/Q1huf8DuAjPOUQ2Se0YZZ4avDa0WadUWeR7W+IZsgHQ5LIct+LR4u1562nhItSoY2ZG
9NRjtBJT/4j/w3cg6uxyCTrZoxL4PEwfr36Yc0zzfTrSxkVJ3fU+4BV7DHDLjX1VWqwdmS79h+vb
gSZ1OveidFrunFNB9xL6A76x/hnkljC85lZG8tt769p5FD4usTwP7HPLjk2CmGqsVqUf/4nFiDQI
93yLQp8DTYnPI+6S5p4E5devyN6yypdiG3jKWZmbXQ9908gPhH6EP/lpiF8F8xt0kmaAhSlvM7ZB
/Lcky0VaZ5qpZo3kfUytWOP5Vo8Yr2B8pfOOSWyiqgwr5zKzXasAXc4+YTHGSF+AXIaTZXCeDjMo
UoU1jXOw5U0oXEn3c2DRLy5jdzbqADYV2ZjJu7xZZlxppv6e6UxQtjV2Hzwj4dD5MdGnHHPHsKGy
Arf4HIwTwme/fg9hwcGv/e+hHd+3Gdr+sqBPlQlcmwfedFjHFxcTaMXPqpkdIZHZIoLDmdiytvLD
l8AmPCSPt8unVfoTdEpmd68EjwEETaQ88VncSRfenzb/hmu9Ln4VRchGZuspxylUqqV8k5UgmxEa
zf4rMLl/o/BJMYYMDL3+CgSsGVvHyGX/rkOgTiVHfHEt5erlD8vFN1ITW9bw2fHs3dHB5kyLT5Rl
62wYIS0zMi6OlSFb/ehDZWcEjqQQO2lD3UuH85g6FuSyzCgykeDV3WHvK4kXxVlirA769e4hNX5p
VeclRxbPTNbDfSlipovBaFrp0ewAec2L3DHcGThQfT0XAeRHEKpQSjnZXR3SOXjpajHspCbivumR
VLBvem44yOqTHqa/ntGGKnF0oDeK8OcuBiruNZ9KROYIJPy0+nnUnQHfF8R3F8DjVgt/YqlyYPBD
aXNc495UuTJT+4gdT7cVQ72/GSbhX+qZsIr12pU0ARtIGIcuMQxZy+syp+UFLf8RTmhZmsPV/JXD
oAHl09fJfKR5PLVxwb/4gnopf5V34N3KRNUjgjIQTY7P1w18PupytmNkSWY7FQyPOmZPvzIOToiC
9zXkLpAi5O94sLZW6CRCPEg1bqaODt7VkJVs8JHQOd3Huj4SkOYMFEZG1i3oy2KFDIgoUXwtGCW2
vXzvaET+vNY8i32QFR9thxyS0D+Al81UGLsJrAnckhoOWJ3lJjDqci8B1I9/fxznIS1EJuZp7StJ
gFAGcKe0P4lC5JghqSN8qY9/Ht2jPaQIbeGM4t9oAaOPS3TlqQzI4uVEe9t3fKvCQQA7x+vH7TAK
6VKyB8UAZ6hUl5uihM/RZTrqEhForui/h7psCbVVKaJV3UtkIFFSUrIHD0h7aePZugWnLV0krk1E
rOE68kFvs47qRG2XvaBNfzR+eG7utPT8O+puOteyGRo/K8bzynF6mX08xsVhKmbNyHkOtTWUTzQv
qBmxdEbmpG2Wj5q9YAPDilyW/VBlXtJX2zzJiU8w0tH9DPeKmOT145wM+gBJdY9CiZI8ctnYJ5SL
inJaxEoQ0Ulq4h6fpg/ESKO+Yj5kSb0oVOYcRHZCXzkpmoiSpVjoYvJkMjh3a053xRgZ0YcQv7s8
C4qCYnls5oYLevXJ9HfKeHRlPOpTmw/2NqkvORJdMJ34JAH3+asPBPgyKxJCaS27UWAAIAbv7G7j
lMkACAHwxYeoXCkGmJ9at+T+TtoYiwk5EfMQa1AjnS4PEcfimHJELp+q4uaCsdMIMvkV9OCL3iQJ
ZRSNM7OvLYZPPSAAMJuIXaG4pQ7G0nIZpVQDInmSg7kBmYXuI1uuED8XQxe7tA/CnfRyg5uXDqLV
DQPwxclzaPsbT1uVqCrXSmCbRd3XmslGGaExshfSn4Km8NczZdnGY09EQBlDXECdkKwYjM2SgSLo
MlEMMLTzC/b9MC5EzDUDjgISBusA6R/aGir5W8nmk8EEjOHN1qb6tS2/nwQiMrVmDX+VPXq/GQrj
U0rTuhjXgViX7Xerr+fSylkc7t25FaSMBIYcSDLdinzl0OFpTm7UMpBFzKUsUUYYyfR0t1gv6HDD
p/cAM1agOS1UvRmOHiS8mxaInTaTiWc5h2ZdfS6fRLIg8kvbn7LNvwCUM6cDUxUKvuZM1PejF7KP
UseyYs6omIEJhN/URZMXmJMEjbFnn8iCn4on3ruasX9QfAxVAT3+YE22V2lj+m+PgrMXI5wHY5Oe
xCiFHgYX9dkBmJWm9CLrmHwKw23AiyLaXTl3Gxj40EzZw7hEEqnnfL6XOEd+j/TDEJyxPA57Eg7K
XkRlvM4/AurjbBO1S4efkpdgUpjEvIQ231ZkBP9lgrWQhvTeG2j1A1oHnBGJ6kBSUqz58mo+pZCz
PN0INnJRXXklQ7YEbd9oK9j9h6IildqN333i8y2DII5XPLeNpcqixmh5mPgHsae+BpUs9r67NlL+
CD/Rn63IKM/A+QX5lSrxRoJ7FfoF2fE8kOB2EPnSFAyGIRJglmVcEhGA5hNtRFM8iEvN759y72t+
Q0qiCcQ/ECFdwu85WDcx52v//bSbqRrjsx1urQWpPvd3D3raUhPmti3Shdg03LIB7J2wEzwDhrMy
m+iR3GolYogcmHGvcli269Kb0jRVBk7trU/VU2VoLaxfIka5geaIlKnbhdI4pUU4EsFalDdM/eS9
BhvOzcWOPaeEwWt72n8DMY7lD+4xL+OiAbOF6lTpFbU5hGA/+wKTSh/N3GVc0/xBshg8KTVb3+W+
aZo4NGu/inDumiYdCcc5Sr3SGPWG6Xc8FCRfleBQ0rHsPDti7mJHc7Kz/Gw3nWsVOvKy0kTpKtXT
Wg9NUMDIcv+YbDQYRfHkkpU5ijERhD4OAlXrmC76QJUfHL2bRIZ3g24V4eBvy15ccE8AhHQcjGqE
XmhjlS7JPqNRVU7S6jsP1LFuQ96mxgeTocOSCNRYz7PD99xHm9wi/vZphYp7sK509DKs6zFL69Dh
bTIgUOpEOR/jGlReBOQmiZfYMK2Hcd6w97WEintCC/IlY+Pt7DY7YASfJmtsNfaHdQrIKKOpH4Vm
YAltFYVyRQNGBUR98vRPjDfKCKYlj2STfdX/et8pFhmtk98Km8WuVqVoQEealRRHzsb3coxRJ3rv
jdxsUQp8fo9srOvswf5uKrWqsW56WwvOs1hV64zRogFNtpcZ10LxE/OAElMFZvnvAKP9eYBk6Y9m
Vns0T3GGZRHqSXLwb3sWPAI+QnGBsQaquXRvioz/JAhP7PPljL6aXUp4vGD5o1tTIEIt2yTyGEON
pdCEhX/GKM4SUHb296COPGBt65jfOZMHvd52KKmsMlJ/7jdk3LF5l3dtyNGWByYRDFPyzof2+Bu/
W3+qPvrXuccmrKefPBE4u6UzASZjYyLiHu6MQVHlfJx6KvUSyxhEz9tpIVGsJUVkQJBDV36Wtyqh
2jmLRtkR54XgAs7Lo5ZYWpxwweEC1ELl42rh/1P9uQ3K/1s9uSVNZE+PCmPXjlY+b8ro/IsFOTk1
nPogVF9rn1oPjyjETzPU3coeVaa7zXuCY7fXj7lHpkSlQevQOcnICcb88SE2UIOE9+sfifvtOjPU
89n3H3ePKM/VPzRTHQSLL4WJU8wBm2bmpsnD8HSDvAAc80VWFLU0AbE5ECeOG/nQC0K9PCS017GK
ejgqQtQuHq5yz+1FcUH0vWGpS1BiZWjbr+LRKz+EE4jVE2586W3FmqDbPwGlijCc7Vwp6g5QHd6u
o5oXnbzrUHKVYpO34qVPBqQRouUOcZJyEzGcDX/R3+eqsNQyRSZMRxsgnKgMCEZMP2qc7f88YiWn
Ls3DjUxCFddPVnFhJmnnWDA+5HO1jN/fI/DVk5+cLsF3GJAKwPhY4Hf6/rmtVBK5kB5aOkk4/ino
Cq7wliZdWYti5aQR/TePwmj2nggxwnzHC0Hy7xTa/E1L/J+lgWNDcKn5qmhlFUdN4lAE+xkYsE53
bPtfWVNDUSuGhgN9eRzbXJ8wM5zygepQx5Hj9xrmHYa9IG0iE2yqIj2qd6ZVlMwsN8/zs/dk8RN/
qtKTdHQINNWxDwDHtHUxbSE1YpUwYjjnLy6JPdoYu3l+x0YDjtU8owEvPLhKLH+2M8pwWVmHrofe
2F7d6BjeqS4z7Xv2fiHgSUNfCF7Fe9FokYjWweD9A3vX2FaO5d+Xw77PMGbYS5jzVPq9gQ6KR2t4
tfWX1jpH8/0scN6NQX9z+Ah04i9HfVpCMI/c3Kqdu9g1ma/YWdJsqLCvMCqtuae4+VtW0xRpFq7i
HLtpAyRs42aA88WrQ2njdoIo3wRHZvJETbZMIwDOf+a4AIChskfo77/t7booVzrre8Mc7fwcONII
2OHRWFwemTr3avhRBwYQrXiJmckCcOB1+Q4E6XVk2N7vp1yrJBGp8AxYM1yDows3KbK1QMHKtacH
yTy0TMCknuKabxz9lLBIVfDiskt/Qh/5OOaUTpiAIYoLyLegpQ/P1iT8yN1c8CkzStZp2haUo+B1
GjBCLF+c3kFfCFgqC8GhOPZvP2cNi0UEwFjCSqHQNN3lYtNoy5nndkwueWdXsK/J/1seoMzuYViI
A1prIhZypQuSRVHcFB4TcZzn4Yf6PbEIEqUxbpBzAqfabCnbSGpIvdbXR8Si/17e/wGeVuZlPYNo
2i1JnE76lv5KNkiJqx6kPmPpOXBx5ys+P89s6VJsOpWOp2Ol6xve4q67YxZ+RhiVIVUU5pix85Tk
JwHNStbmmc1CD7nmYxq1vfnjoO/G+snK/NlvBAfsaZaD/2bpw1uS1BeATH9YqlcZ9vo+EGH4VnKI
A3ge027iC6f8QXPZRzfSgk3Ax87AkGCutX0bH44LS8+JZcmPS3373jzfOTDJHaEE36G7aBYkKGCl
1LZcoaebfBrlHLwK6+6OH7cMFp3noYFfgk0tjdAVxx1O/mO6btT9Q2eqOeQj3tPFqCZZIpuj91kx
iaSOJITTYdih+Hc8EGQNMh4IOtj59MT0Jt6Z0xj2t71iVCf67mnZwqyErqV3sdrkNnxqKU3t/FFi
4aJ56J9cYxOrABVHQoWOk6nuLokbvcF/RSEyTl/k+fynFk4omwmwda5bYvc13QOGrZ+bngJzkHQa
+XVf4nbUZsgLgVtTiyMuZYR6ZsnNOCDTI3I4nw6EXJG9w16q6gtfHcwpO8jkbxEkaSqbgLLrqSTJ
gQU6sDrab4Le57CtGyJXbu0Z3q7kNswIs/2bieLUE9ZQi6V4/+bJ+pmQ+5fziSFwnjwr1MEdINtB
dKaSFkNADZUjdvcR7RXqTspHaIAkqWS4pparDGREOMKaM95TzAPNHTcYnFAJHNSjSG2O45Gv/Kdw
+dtTyqupF+QPx19ismLisPqlw6Mn0qcQOqQFs8D5lLdrD+Og1KbMjQ6Kcy82kK4xtHtuCl5bmLlb
CUj3id+dTNxHbv0LHe34qruZF+HtvkS/zKqI+xP1tg31LuLI5ePvzNbOfMIz+TJECMRvLuXuRY00
3ot7ruNFOOLSP/uR8f/utaDzir4WyV/4ioPGkxZgu530lkw4WlJ26Xh+5xSf2NOTFGaInVoGoNgq
GIkbOTJoupQtAqe6qf/RkZJQyv9Dty6MW74Rio2JjR6d/lUn51J/XSdkbnhXAOTh4nAarJOYm8v4
MPA+HhR+VacZxIQbj3JFn+Z0t/rKJCKwutikWwOuWcXPAvp4KRa6P/VdkqHxVwoKK3h/8nr26UOv
LOAu+ZPJSbX2PITVYyEqv5QPoovUr7RWKsmij0KO4Ylp5/QFgz9GVYDaEYpoGVlKNrgZxJffkwTS
ok6VM3n6QGDYksSYvRrHBmUcCoEHDlk0Az2GDnrq7BQQ9NwzdqCJIHqiVj5YH3TsDryUXZWCqkmV
vZF6LZv/0pBfZS0RCsZfMIy1gHcvWxGUQTFWfJD/duMWE0ggkMw24RRp2yxe5eGaTWosXfVWqMJC
eTfttGQeoK1pfd344Kn+Fw/AubZ6u0nSiD80TiEbM9z4/NkTKxeN8iwrNrw6GadvcSg5JtK+n+n/
PLLB8exH0M13Nw6W78XSePLjdl+FBstfOV9Az5VBWRM/SokaViCoEwgIuuzqoQAm7WCwVGQj4VpA
uG6gRyNnT8uMegzV/TmJyaRLWVXP5JCcPPj7wqlVSJGKG2RX53E5BFzaevYJlZcSxpi2cp83G27J
sbkKFBcPjtmezOPTxILnb/mm4XsUeKyphO3wR150WLnf1iZ2PXqJzvUt0jo8aYY5QMtwoD3tkQ3m
7F4GLyEaFEnZ6STdJEKEYULZoMPBiBa1jVpWOCAwSIop+8QAXDTMWcnO8GY6R4hyMozascBPb2xL
lBf4ZiSDem84yBpZ2/UdwWb2ZzyF5WvLZiE7Zly5/Grb7kA/dolYrf3xH4Pk8a2i4faQNH8Ek49n
TqOnC/OHDWJpizptEnUBNqJt4ZJX/emOQkVPRYPMy14a/c/h8C70bMmax1njMPBuklyRezy6Hm2e
PMGYMZOYOnQgii3aficfSXAI0pKx75lJ9EG9DZfHGYGPwTTTdUCankwjtIOCGb23E+Wgw/eaI3uP
zQ1P1j2I67uo34E/utUaPPpNt+EmwesvsZvcQ4JH7i9Jw5Gr+Xg47VFK0Dwsm2CPyWzLsKR+p2bm
mBaK0p1JIXu5v4X0qFtSqdE6hZCXYw6dfTYx/vNnINUZSvZGBAW4SGckFWeVOd0SLRqndg5Oa0aC
8dcazNqp5Tt/R0iG4glmM9VP7a1R5NbtDS1+XNQdl7BH93j4p3EBzROjrzC0cywnGwBxFkubpmWW
jC4XHHI9RLFcD+Cbp+JHTAbL+DnVRtxCU3a2JUOV48M+iuHLEY/GrTOIG27+J5nYm7Z6JUx8EgQL
THaCmw15HGi59QDGsZSM7JdwQ9DTR0gTfOXmgIYrZVUoJVZ6QYmPLkqTT0CZpglzgG4KCHJGtxD8
VDfWybnylT5XzH+5L9Y3ODKcqd6k6KEVzhWlL9E87kwDBHZjrVUlLQEbvy6ApY+yNvCzQBIXIZr6
BxEBrAThaIqJX5BQ1HRCieohgLBZwhieytP1gexPrnN+tqKAYs4yvvo04FwvfEEyalqz1G2doKn+
UlTitDoSfR58qZS20ptdCiMPhjr7bdjv0VQfOlubYq6rAKgNpXg1TRzDPU8wnSLQ0ydVaMy84/c7
2evALGklE7TI0apmrz0pBh3xRFh4wVZTlhNbyC3tYesOWjklFU0wbUoxViihpyiPPaXJnv7F9mAy
ZdTGntEVU6OzS8dZonOqfcGM8dofTJNsAbEtrVSCTJsC1gQNDF52QT8PoKz16VQHYk6GM0cWKxDR
nzi0VRImMghdFW2kH8nNPnuY3l/EiPM8WkG+9DeRsxr1uXdldXUtY7Ik4UUI1t4AX/o/FQkOfsgX
yoRCV7sm5jw7oowHs03Yr0R2vJYXsZGhKaC+D2YPOwWik3iV0QW4eOy/L02m4ZwKERDz1LQbcuJ7
bHg+0Pzco4vHLgvR/i/Sf1wMAoyEbUAChWfMQPZSzG0wnTE3Kn5Evuq/YbOPXLfMaD8VS92ey8Zd
EFkdPh2CE7Mc4Api79qu2RsHNIqOPx4Nc8U8dff78as/ZfxVEltOin9a8camZqgiR3G6Vlb93bjl
JlZtYiXobOm+kTIlpe8fHVQSUeJj0sO5Fg0hGVF7Acefvxy2RzH2KRQ9l0xigTqP9pzYpSPd6Jut
iEKiw/u9JvZo/mMMXaDHHK6OKFIqk9bfYcD02J0y0WZ3edDXXG+ltP7WzjSWXBun2IFWaI1JPbz1
OHhXcm5bK0RCZ0rDQupNYIDm5Lu+rO83Pwdsj8JQxnsYDnB3KsJDoA2LqMEY2brlRMGN6zc6wSj+
sgsTr3T2O+86GUtNJcj5aMgcFFJfAtcDXLMrSKxI28wq2epuLcUuAHMV6ZapnAjmu8o+ctlQMgot
xYYZYnv7bHJePJeqOvxz+4WYx2/ZfMMQZXhzfFjOSTD5XiDoVWW101q1vlJb4FjJmrOfVKxWL+Kb
z7P88TewAeO7feqvlehd7+XFQvYx1+4qBmcWJkZvmpXH5sFUdiJcIDAVb9Fa1sNeJZutf66YGAHi
8VJE171yJVQ9kLCA3M6WFE7ffb26dWK+Xjs0YyVZkzt+UjDNgvFjjN72qgjgOv+Ay7tZoxu0jGGL
KHoQ0gefGjTT1pZSnXUVyB3JxHjt5RF/hIshJCVVcV198lFUgIks2ng/NtM3EI6CiZ27AT1WRayP
KNUsMkFBBL36LLRSw8OYFMODYEjsElWtoIjhNcOJ+33hIUGa+7JHIQ3kHBtF9gi6fwosxBwAnIZ4
Ot7v2gCgCP8G5brHMkkFoRPdKFE8Cc0gsNT2ZGA+c9V7k98bZmzJV+fA0u5lFRwOsm5cuCtxdYpC
6prJpjnLD074tNqkRHwEjs4GpRkNmZZg4NGPK3ooY5PbVhg2jfKaAkz7f+DHa/XtFkjdbLXAwcfY
/u7uGn+qGbZktRCXeaghXJ7vOzXaRmd/m27f0dibjiM9Hd2uNPk4dKFUU2OGkY5xNMtj+w4+LpQH
86NEmPw/QFN1vdBpiS4+nEwML6J6N8BvG1H9OReI2RtQ+CKwrRA+shn/R6vmcwIZ7dE6Lb3ggGfz
ikT0uEoCPhvxFsXm3pQSvj4vM7F+8zgTVhOR2nRlopZ+ET8MWmjP54EnW29Rn3T4cFwYQJH3Be8i
FfTQ7Som7tdxxgkkV2XeL9NfAG9m79ZgGEhsaREAWzjzvukksAUjcVLsAvBt0VmY9vJRzrz+sw4B
Bn01p6u/qcgTF0f84+wLTDiHxtwT/FpD3JWdpfPFGbBHkHFM/0OwT0dhAcgqriNVs3TisBCa/TRY
fAUWuYL2QaRDEQ7zvz5qlMQWWV2VoHWUVyBaqVvFAwY+yt54ygLMbqi1ipXikeet2NkTsOFuqH7s
3+yJkp8SDxKByGPAJd/gsSQPCHX0RXHaWe8YfR451VetgseP/3rQE6PI34+kZ2ZP0icf5KkEXlQ+
JfQQJe9hfxTJAkcny+RnkYTSrIgMrhQwAZ46+Dfu0VFmnGwjE7/KitEEJQnRr5b6wSJzlZXY1FO2
t8RLOeWm2aTkAj9Kl2PaG18WxTsLfQhQhQ+ARNLVb3egi3glk1myTfteRUzyJFDFOUu/kXQiUr10
7dLB7UVA80uNaal4MxTL8FBQkR9Bjz7DGurs3l7xCAiVD1XgGAp4uk7Z4UTe/9GyEzJXTTiM+Tmf
ZAHSb7HDTWs5s5V04xLUi17M2wEFg38vfptRyoIcR+nCKBwm7Ff72RP5sIMjXF3g0By8eTe2vqYG
xe0VCN8Z00GZFDZi53kXa512oTjEjT/2kOlSgKwSs9IVrUiIrzD5zFVvyKq2F9qgOf9Gepa9T2d7
Yhb1ZshWuKOwjwF1/cgJosj5PUUC9YH0PgEzVnbaeJzoUg31wc/WcD5TMXvQNDemHeT8szg+CAkY
MZQpxEgnmf3f/OA9q6wTG4Okv22OgCMMEKLc18hIP0rO9eUAXBYkSjFhl0XJFaRxvwrulk6cJMYF
hduSCyLkfNNVJ9U2xOqe2Yj39/gAe5T5E5rAl/Uonp3A3rK3GavAxgpaowrWdJN6mxr3qUYB8Ie2
+eU1Nm9hVoKqbuBVYDqcr2YOTkFO8gwCFN/TB7Cw1GyHGi3EH7XYG78gavSLwNdV2XFVBDMtzvu0
kn/w/BSWorFAFiHo+VKMBD1On1Oew69MZAnGzqsFORusxLXMAxiHyBnKfPzn+tu6CwbKBietAbbG
2SKGcG+DK5ig+vRMYRojZwmCzRsF0ecnqzqp2VeXf/TDjMW1rIbWeSkG/7QxOpAThOp29KjCREK7
QtD6+g9XJSj7BdUti0ZqYAX0nfhRADVRLeYUtUfdKNqD4Ngo0bKdJo4pB86f4r4Lh24JkDIKfNzh
gEA2PzPjWSXDvXkKJyc4vo6tf85jOk6UYBkg1IlJO1J8eUYXNCtNNqezGff/rlOR/7w0AUGn+8x5
yJOg348OdnmILokULnSUP1MS8w5zvJQ5rvma71mUY7OpCv+kSpp9NpWkBuTuzfxSKrgl+9txWLTX
9M4SI36Tmh6bukeKJwmQ9myPBOX3HH4WAz+lAfbN2akodKC7JeY+LyU7gKJXLgHYOlhsNfSNeoiF
DGvxcjpuY4EI3/h+LvyRNFIA6cGPturvBX86Foo2mUXgAYAlUO5jj7ky32q7+ZcpKTyrbwjh0Wqc
/9SYwCadDZ7YG6xRuMUcLLpjRArMTeRf+yXfQV0O3Z0/mnCUpx33Dvr7ISqZYe6mNs3uy/XZ1WGd
1RnGmQT2Whtr3eTfOhdUxYVr1V/Vrm3o4QXfo++iSF/Ij4vR9s/yY1ue2fKRf+/Wvs9YXxYwaI5i
GEHw+nhTilkJ1Qbap4cdKP0ZavjqPzaxGiIljO1YLh2IwSvCc2QkxnySN44NaF0eJiLT+k1Z5/EE
cyrg3hBY8QK6e7DTG5XI459RnSsvhfXuxBh9JEbbttOOi1YwjM/Najo0yEhtlcaGBiMmC2ybaznb
R8+WjQdnqklcNSJ887i5skYdcDWkFIIurEeMbo7bo3U8Qi8xLohyw0o5u2wy1/sebvDrjkymfGNe
Bj+1Iyks9sD4dTY0UFHRb7j6WCaDQdQrCD5GnffjeyTNjGlcvAVsoXCpw82wYGRjr6I+3Uzz+An4
sVwyA7drFb2VFLvO1hixRDwkPbifQSxnufQF4N+KscCX+yvDWc/zezctyt0KqAGDwGlioZCUVe16
4/6R54fuYQux4tDJgF6P8An5W37FADJ1Ia6dfRC6/zNWejbSE3iT2/+dfRFKnVWdxh56I7wceKOc
oWxL8GM9m/WGR5T7mLUbxwuJZXK0f11+jdny+7OppaLjbqeorqZFaylDGF+1ZDDZUrnMlg8hSVj5
PtyShrPQf4rCgQGA3u4ZXmWMzKa86Ju/qrRCp/SYYyCuyjuPvchZQVMuOjY+LzH3QUvNJD3n67XQ
FtahrLotC5La5ITuTSgBxvbnmWBZaJBSB9DOuGFU7QVY8MAr25nIOsHJ5+w85QS0h2CkZJMr1tJN
BMRKgYPMs/30TvDym93CO5GLuCsAFOuiSDdollkCYn+3GwZa0ZFPeNzX1Zx6qUESoyEapdF7KCv9
gtTWwS4QQaggAeW6Cnfj2yIfQkHwfbnsSHemj37doZB1K98D7VW19MRgXSD/lmlSxquxMlIK7Iy/
I5DHTiupAIQbfH9HmMNeh0b9r0jQ09r/Fw+/xAw0dyenYzEKEAEcBjkLBp7+Jzk7o8EF89ylBPgG
WAaAHJIyH6M6BHE6z5O88XPecqhhhyKsilyh21gi3YirImx6OGaEtyR+XV5ObPxSDXQ1SjFsYltS
mmcs50IT9SrG0l2lcI1k9oalTCRFD95Q75hfghWpBWqCu8Lb3YyzKa+3FRl+n4MFJWtzzZTsA7nd
E+yMGq6TfeWNjYep3FtXiyi6N+XBjcG6FaV/+sqviy1f/JmYFul+O+oqU0mFBhqpdFCq9kaW7tmi
8YV1AmAfEEypdPuI8ndYoobqESa5WamXrglhB7UqLP1gSRkDWrx4waVCc+4fa3m6qyWN/tyKi5MC
B7N68ad5omF8HG4vI9eBMQQ6+aRarxBK1u1Gu6xps+dUvXM11a9f8ZjSPyessDkvYaTXyhAq4N9D
B3eg4SwNIMybz2dyNoDAPk/pssv3ySdKk5FFq3fZnp+F7TzYrKAtLKtXlOpqNB0ApSDvvXutP9xk
6N8eoCf5U5d7NFR8Zx9BJcfLnqRE/oe4WE4yNJoB4XjhBnT7+x87GsAJ7dD9Tams+4sht8z/EiSq
wtoJmfMxEpmTSoJtaqi6FGNHfqxbmtDuDCmM29lm2nxH36XhHH/Ga8BLCKyP8XKxwXwj1Lum+Jkp
Poq3VTMgqd+2KEasnfeDbe13HqY+2skoVRO/VO3GxWnnIRO0KfCAMsPuBAA1aNfdJCS2/vvU56Xr
XE9hqyGy7QUi1pQ2j+ivjJs8VCr32XXgESgvCFc1B6aQGgUQTOd9m1KLxO98qyrwYc+POXwADLmX
pN3EXMihyGj+Q399UVvKWoiu0IPngsZHIC37G5+LxrZm27nfLXSC7iRVkizU9noFFwbjkQ2OM4jy
kLKgbrnFZpi1teUqx0wsue4y5ihN5sfnICIjWccAskfFoVXe5+l9+l+Aa48IRSgo/0uKvRHKrQOD
pMRRUK44HAHTYOfXADpfeQ5EmldmWjHQUF9uB4/Ns32tcOmnHk5G+fXofAXzMyspviPFMDx4OL7h
ssZ9NAz1u9EGskofRtjXtfy/cGOvONGOFB+/4K9X9D/VYaMZoxhVQ5p7xFf8gKnwC2UZDIQFcAq5
Ur93lmHuuYDY133g/8hudxk6oTFRS4wQNbmuh/gRqV47RvxbEa2jxs2ij0Ta04FZmLVuQeyhAn6c
aB/aQauU3RfOYMGMR0APBw4S9BR529VVFZwOS4kelEoAiINNN0JS5LrkOPp5z+FaCB1IPOsRRb6X
dFAx7ckMasvZQgqUM5hbxi8o8I6Hzg2bq+flG8PuD9JI54QA+DWKUVLVnbYe4UsEaJ0Qv8rYZjRu
7itrBctcqr095wPNcVkq3rg9CEm2RlLchzQzPFh6rKK8V7gxWqW7CThqRAn+oHKJxYdUKmhhTRao
tFiNYbzOvTELRXMKdZPNR9Fgp/S806ypInYFgt92UitKVZkaLsEDsV5CT/CR7rDURDv6qK1r/FJv
WC7NbqV9/LDCybvl8llm10Q+Jh2Rqb+jUpCLykMvAGNqj+D4YPh/J9rX4EKXzTh6Fw94060XQn++
jIcVcz4ciUwrjXgZhebl6sXM5tM3lX44CDJzRe31eBsFWlrL0eDalg9l2B/ZFTsBFv4YK0M2V7hk
zq25wgL3npQj1382I7SZ88+vCVyakOPQkBeLiMHUUs/8F4BcQLgHoW3I6O6eNQQ7x+cpCEr/2hEx
jDdO8e4MYtryjw2WZKKwUOTU5AzjvIzmjGeYgYWTZnSig98yNeJWtIAAQ48fDjLjsDS1P3ahwceQ
IEsfG0vaLTU4ml87m4gpW0X27dRdC53Cm5p8TA29NSYkwkUIWN483wuR65I6A+2s6Pkau0FwHB7j
DFaQb7VudP3tpWOnDvbteE0QNzxso6RUUvk4J3zYiqUdjO92NegE6P2bOUmUcNrgI+mAtvxd+Ihn
A+Wb4VuRgJolcByAARK2xbt6j+BtR33NijMz4ucoA9wH6yPFRQZxWcL1p6csIQbReiM4beb4Jgkd
mGdc5ncbKxT6LAnKu/7AKMzDmSOY6qZhm1rmc38kyI3+d5qWDslawuJdczzB4BRjSUrQkO+44HTq
eysq47qLN5BdpskQwEdp/94S3yMhAr1poIj3KZlh88OQN1dObpeYeMJEgNuwVrHFD2qmfDdbiCjk
bGZBpyuVge2K5tmc/fHse2xrmRKgRBgwogibySzLUOpkVFJkFNT/nkmDOZD3wpSBlXp8aI6k+GMx
IH94Sjj3mpLjS5X/4knm3hXMXadN6m+SCS8cuR6SiRIvI2Cw5L4UfE/jfuXMnxWRheXVW9LCTN2T
FnZQPlQcCts1GRwJ+IpjceICaeHxbBrftwcD36IdrukilRKS9edcSqGfkNuihAEXrpfDTZjN89Jh
Wx07OuY0yZiH5XnwV0sJpqNy/PzLdhUVS+zIz4ahiMG5dkHhxMurTeTeMdqMzmgvspCtrxOwsPUp
zGfN9vWmPWoqilPcKgN0Wgy9FhyNuqKRM6aqeZejiRAwTGTiAx+q5d/JoMFiRFM/yBUKyLvlWzbQ
TE0DtHsJagMXjIOp2r81I11eFedMWGVlSkGiAAG8cdkhJ7TE65Wk8+304ryjhmKihotU8M6/VjqY
1lyHhAF3QeLLc31kvel45n/RRdBtC/a84Z8iqAILoubD8y+8KmJ3dIQsu+NoIg9rAUrtkZiU+WQp
97PN/shoh1BiJlHSzzKZfU63HzBzkXyRlaHHoNuQ+rvcK2uGB51e8PMFJynuJreuvslEAcBTI2GV
AZOWvi0pj9W2K5+1Hy6R3E6jtQsd3Q+OhU1hQaHXuDpEqKE/NCHgIBUNZMgj6o9ADiHa7ZBWkZJx
wIO6C6owG0YGJtHEdQuL6PmYu/zzmb6bgMUH6NyONzKi2vhnqVw8dkAjmVTL7lF6mPdkMgdiLnbf
HQYPmlf8/HM5PBBozA1KI3t9gtDEiByNDp7i/tTuiV+oOI/nNsuVY7WppeiYcMOg+H7Q+8dATivU
CuEniCN3k/Xdhh3q/XSMU3fpjBZ0QAKbVgrmGSUofp44VjHRF19opvfVl6Cge38L7toVZvuN76bn
RZxKjFoTILv544OwvOhfOPhF07YQvRcWw3vjo5rgyF1wHJ7uKd1WPKBKfgT4hDh1y8SbOqUBeDgM
ckeDFTeRDdWmBdr76DE3VF8mCzwQgzGir9ZVi1gp187NXLpBsa/4M0dY3NdLU4kTjCNhcJRvJlE2
qdNMIHugqQEtpLFbz9+pT2zULCsryp5BbS9p2rIkpyj7oa5WZEXoQ6Qk1KRfiqpsHWjB2D6hPOhQ
kI6KxBJE8FOKXWD1qFQ+ktm3D6X9XyHFtvq+GWkbtu+YVkpZOEI/l9D1L00FKWmL/IsWeAKyOn/m
b81jHdT89ZYmz76941CqPp6n+jS4aJSzcS9VtIVTuNhN50yYsJ92bbu9uoFdMXMAMswv33U08lxH
J6qHxtHWnigE7Q0Ro1GWjN2mx5FLQFLBXPeg24LuSH7uCIVi07a2cKic44bfChOlbTR9/IgbrqQe
Oq4b73C5q7/4B2p1CuZnzpDAL5ulnQmbrmIzITbwZ2PcL1wifs38YbpNJPLpHpepbUYRhnYhESxz
94gBsyePWSOdhSR0no7qoDnvMiUZGGo4/uarWB5Ob1aElKzoxM0O1Tp+4psjqryZdGJ28Kne7I1V
jro50epkyfK0675Rkpd0wy/LB1wAITSVQIL3+esz154KMvQB5/IyjzOV/1zVKhcvIuylTz03SUYK
mzEZxJmPQhLaJ9CFhCsqyrEMAj2p2RtLSYwd7ZBFdS+q/Md5XYLWHbSx7//q1jp7Eg1KqoSfq/Gp
JhCYP04cL5Pskn0cSq/fHjPxAKm6QinuJ7bwyITFl0YdS8o835xbaYMieS54FzQHpY4sbSKFZhmA
BI6cpM5F3GHPT+ZhhJ7g7BB7dSJnos+L8x1dAkXLBukrMu9zs6uvScJOJ8xVJ1+0mTTtFe29bOV8
i6Ed2ql9Z2ER5V8KKakuaYLLwR60Y3FF4BUytslddgKOOWCiZAelh3c+pxY7VvomlbqEZrau4ASP
vb8FHTU1cu//b3u2kfA/WWswU3yaZ1jcEAo4q34ILdbQ9arTHp8MDt9iX8y2zJsvfqIv2y1o02BQ
w8ObWNyPG/bhe5l6rarc6Kk4ZRsbCHeCX2VsQkHgzMxBAykLXqYDRuK77U1JiRd/TxiKuW+3ld4A
3H7do7JxbD2gywAa9r/I1DoaA3D0YrSydaFEjPdp36+da9hC2Oh7Vef9UL+vQs7TwsG8rC0w7bDk
l3cJUh55+WBNaewictsEPiUn8mh/s4XB0/tcz9MUzK4W06w9ppPNW/lPaBJuZrzp0bCgXT0Vi35O
vEfZSwU+RCF7wuE4RyVp3QyP46aiP9mGnFQYRMMtVkiBUDp8Ya8e7v7rKpzmwOU/x2aOxAi41MSc
PsHrS+nlrjW7f8T8TXzRqJov/TMo+z5sPM6zVQh+imK7/EJVGDIJT+cfSRFbfvcRBLRJpiBGdztn
05SBE5YRGC/jIJoINIX9+r55sFyKmmCUn/s2nCI3grz6BgQ/ymntdBR8FEdYEQd1lHyd3v76/r/L
ftz7SiZirQXSJQ2dBpcqu8UkZ4mDCIn8bcvzhDNEUCqfvTdgO7gNPKpzQmTJzgNUI6vM0SrgYE6s
eGipeXE5UDqFiZje7lFwPM9Da4kM+G43jmBvOcvRsmo9h7R0/ereU5el3uPicvD4ujlcIcUQAYXc
FxLx8KsNBuwhmTQG7i00fq3NS9r8iOKytuUajJtJY+6RdNE+e5R3HS4JY1CjQSM3GxJ3OqWgeEzf
4a13qc93BhraMl7P+mdjNlkFwTl579P268sJWUMJ5uNaD5br4DCcmmLGdzl5iIK2DXFvETtWAghp
1KEXTRNzkITmlE8QXtynec/4gvFPCxAGoAa3V7yyhkkyWj2xwnXgH95cfswgzK+M/8CGJ+KeI18p
z132B0RdWjkQcjJPzpc5dPDT8Lii68d6mxoMOkP6JEyRdfPgsCD5aDs2O1w4RU5L1V+LRMT2YSls
A+T58zWxH9lXS7uL2MpH2eUshN/rLiA9DvgRi4UfhgORZPnP3mYvuawnlie8kRBZUNQBhlmKVgHR
nBNpA/DEYdXMQyynKt5jhsRYvIzXZq4g3IS+5PmY6vIDOpLGrBFLAVGZ3RH6LdBmm5boD0woAFtV
3FuiibpQKY1ZEx0F7ovgOixBdDeNi1L1AhDueHEPXvaRMvpQ7gW0/GCv+XkzAihUbbKlE0Psa4qz
fw3tnwQWlrwiIsDSQo+JCVtiD3vv9rS9E7GXcwxi2WgMCefSPLM6j1K+t8YBQYZsbb4JwhuO0OF7
AZLjDHiFnqRc9EYYHDNfS3chJSJWHw8mOu4otXjpbJ/vLykmAjvHLV3HNcmtb0eiKFh1rV5YeHvG
gSMD32U8eanWIrkvN9c4HNmEN9WmGa6+tfc//VPuaMA6fIAnFcj/WuUrGFa3j8lNwh3TxfYP4+Zf
tOwoGlnD/BaVVEOMA4BprUwTPqSM1Q55IGltWOz+me821DaK7X49e1qQCAJ7M7qrevxZ3D0aE8EY
wxATNyXEDBPS1MJFCvjqrCDIAS46gQTQKyBCHu0TOeSXwMYCxE0lTQJJU6wGTZNPxb39lMGBXKsa
3sZyVwJ1/gQsCUd9WmC4/qjWbR39DMutPh5ts9u3krSX6c4qjTy1NvZDsdFIX35sqm1Fb4R0QVx7
ID0MMJOG9y5JdHM64Swk1FKQSE4z1+/dh95ls4qXw2KEl4eHmexNlYonwSPcDID1aWXwjqikEyw4
NYNztK8HLjsYiO3FnjlqWHn3WPkcyXERSZfBJ472dxXMPuX07SWVGPPsRBFbn7aTr54NMfXQZQaN
3CND4Jfj+Tlfc6kFLF/8kjfjALJygNf97yFD+NcCpc3oTuV9DvTCWql4acKY4gqsq1wC7CZlAPIO
jBoXcIAcxMUFAWbP4Vr9LEjVoyZETG7ZylyPNo9Nd9A3avbHNJqzh5A5VG30Lp882zWP3hRqKlME
yu7QsazHL6QWnxVlh6/QlJPLgwtL2hxBrGlf654Eh6BzAFvqkFuyN0iNPDyEB76wr7XGqYIk/Yzs
2ENHYa11/qo+czOl5Co3kNAbN19ZOyuhWlcOAjZbxzaUEkYf3CPAzDHS9jDYJnWYwrnwSgDTVcgw
AajuJjdvBoLhhVrvi3+kTJFzWnM0IMgQ8lrje6RxyGkYAB6QUYtv3fe93jP3wPXJdB1Zs1cSimLy
oFoRJqUCBnQJx9pH5fklOz9C+e84TayFLxSMwLQ12YFyScTJK8A2LVFPMwEFS5DacLKhuW8b3YSJ
GfgTXVin4yw6co1XMkI3yI81Wmr16KjVpmspqlwolK7j6MYBOffzhctQf6U0XFk1UJ5/qlOQ1gAm
X57Jc7gkK3cfkbDiq4DccLyLrFbNx38DlubzyLAyeDjhs6ooYEQmto93sWLgA4oK4+8vGtuhgDhf
COBgQJjHIU1WymY9Z2DN7wnBLwLIQkICMLJqLDZFQXkjfgPUwi6x3emnHPR7HGTIvlpm6w9zxTI5
jPFHUif0qLamY7jm5tbzuI1HoCCpwd+MerUhLF7fGhmep7U6PaQp+8OqiV4StOZ4aDc7fp/WHOtf
kw6MB7WPipaPtze80mB5aW37yo2JWXT7XrP6chtJlKZzT3eGXiLICfzPPIcS3v/huqSRvr4FRKbN
W7y7wrQtWe/gppBMRNCbXMuEz+LVu45jSAQGhyzW/CoAyp0RZXrLbtC5moPhH2vLHfMNgvPd0suy
nRKR12cVYEDjGLE70pJr+8WOtbnJFNxw51eZ8KQpoovz8C/r0tbNEujUlfDyvnmYgUx4CNLU4C1q
80A7kuRwNVaPXqNKMGEnOZeCsvIkXLCPtK1vKzvbTDjVUycbZe10Y/LHYdcECyDOqviWxGOv2D7H
Xw4rAuhh0pqspeVpURIobMNOGg3YvetxVjP2t7Xu8pYBpjn/1ZuPJPNudAEXt3nCpYwPWg+CxbIp
3N9g9IpuXF3L1bMLV7CTV+Fp2e/+N4lhePsScCePUgn5LY83bIs6ExDRlYMg8bR/3YC7ZrYdZvNE
emcR/8rQrhyHerbyIH8FrKVnOOtdVPBiBxrlQww84kgCu3V/zQMrtYy9rSevH7hHH6nEL4VE1sO8
wGUeqTWgMncnoQeDLd1BiNT9Nio+IkaHzVK06k8bWUM+2hlmU1SBSWuosf4IRkI/ICMy+KaK4O5h
Hqi2yC/pVASAJVCvPlPIclXInN/eGRic/Tgqz6fWi3yqHrOvWuhFTlzov2X6vioFoTck9A85z/LM
ctuTSa6rXNpdznAO3yVevjzirtTooEuX7ANKhKAD7/BGEgo0wUjpbSVlSp5+diR/JtRhGKDBmy5j
ZkJpWRX0atSDYStwrD/I+IRnFtxbDI11EHvWb/JEbwSsVofVb0s4m9Z5G9qGOyY5hQeQsVZwQpkZ
3mJAIHk0I8qksXvvw1K8cDZa3XT9DT40cX3IOBGtmz86opnIzLvDvKUpcik3BiNgR0MedYDc8GwD
Tyj5pL83IYEH6+Z6klVNrObJ2HP22nDvGRzqOQCBvYZ2sAC9ZfLyS1C2Ur8g9EZF9mheQWCYz3F4
1gkTl4sftGdsw7FksDnvXLp6hAOAQP1JJqJ7ST9/YloZEI93VNRSIm39g8+xyRwWhd3wS+nO+MDR
d89GA5tKNrRk78HHXQdBOyz1eN4lbgbP9VRaCpDt0mKavaRAC+GtnpgRWDG3QTi62hUalee6+VMn
YZtwHT6LPbhtQPULpwE6BpgKpvgkW+zdtQc/4DUqorrXez/JaXUj5nWMRasY2Kas/yBH0J64QPvL
OYLumZlU1oiDHSWPibvkfd+M6f7tB3xp30/sbU6PwhEYNldj/9d3G7KhMHFpX3iafIp5AZuKC5uz
EdAqcccoQrCadxE5wfo0Mhfi/+HSKAdPXAnzV2zFrl2gtXxn2A4dEyfTxW0H0puMSLdklpE6pZIa
2eZWhnazYHlLIqlbmzTA7nYWbplDmH3a9ZQ0xBJ0VbmyX+5MYSqatmD8YP0sSn952H2czhW5R0Bv
vA3JY4ilaVdeykJRxmqwivz65HYnkjtMtqJzQHgfozQexJ95ywVtuSXCzTNP+wZGQjQu+sjhV1rQ
D5q1sbLBn2eg6WvesAuv4EPL6DEcAMuSwVqT7J2x1WE0WH2HrKdqsjo+du01clw6PnoTC+T+Xp3X
ccg3JQ3r9eHvVpChTav4bSxaZlfMFwFuc9tzgCWFOzHtsSjbQn7Iv6Ma7Hy0mEXO9tUonJk4P4dO
YT8YY5mrotVCnZf8wYkSVlMymgzMclUWyfEfmmogg8b96f4ZwDz4lRlSyJW7bAZa5Y81DIEBHzqD
6sUnHYbmxOOGy2vMA0olpS4bwMbypnWH3CA/thArU0wJhQlAEFhUCs+0Wk+rbjqZIsexW4IBos1X
7p8cGHguTzjfOEUdRxcVpwAisAzfCGA5bey++37sfuUj3D9yc5pQAmU41fO+0Djc3SCdlYU3okbd
puZiXdiiqzxmPE0IEs0ns0RLIXtUr+34RnhWMyNZmmP9otnvTEYp8ZOGQzR/w8GspPTpAcJs12dH
owOXVvOZOcK9R0j8RemXU9fghwRizk1xjvvoU4YZ1ONJ7y5kGX2J3B9kJCslmXIyNMMXBg4bd2I4
vth2mBWcMPHlo7uYQwW2355RJw3eOwyYUYJetJ4f3ZyVkOp9sHZPpe9O9+W1X8aZbd+VWc+r7Gx4
Ce89Frz1g9qSsaZpa2KaRGumAVRCRgsnSYyxNe/W+e/yOa3szPT/CF+pJj/xKneBSXgQUwfbsIBU
mUgG28ko3SLmUFStpVdN3VQO+tciXTHopGXHIWG0ocS1A73tnFU8lAQ1T6BsBo5n0xEH4OdRxeCD
LvGfwMb1LhBgoOVgByuc1wh52sdMhI2j5sMoHLb/P1zXgRSLOIKkSmtZL4UeAgHq8U8345/w14Tc
pOswqCypQcQtAA9HDnfCvActXk4KDRxu3av+hDBHquGC26OFaUVInbCyoNidufDnKEjXXK3wHMIg
/C/1EtIoQRyvaNNbIkbD/t5tK0nWefHeaFXzOD50QT2u9QuRWihUoU3dO8Tci+4Y7b6iUftv+N7r
lPri5na6x12GDPJPbJtPk7MUh4K5Hi4liNMCHgeepSyFoIcm3n21oqGE6/Hnci62iZfh58C4yZvd
m5IR49UbKaEahQxNokxUwiCgfhsOmCJUXW9ON3yDOBX7bh0mA1gklbQH5SIqnC2LOi4/cjE/YhX/
n9HkBhVFS5JM0W+jES6Dr2cNZEcKMAxM2QTAQOWm9nW1YkYWrbDOCqXE4rC3SW6CoTjNs8ETT0Dq
G0Nz9MGzhaTZcFkt4m21A32nY5EI43w38jO6q6nFhYTQRz5ypBW3yqJzqHCX0Usgnpt2i9fVeS4x
HGVCR9zbgIHfvWJyjatq/7wjTaiBd+Hn8GRzFXcQBRgj3nIjfWbPEmsZZFDwEAjwLG7omuiTOgoE
2QDU91/C2PspYfkCNSqDJELWuzno3df0AoCicX50i4VgdNaOL+5MdswYhltla1ubIIHX9Oxi/ZYF
o4kyQuXlFqNhA9PHuz2qva7KfNb6DL1t2WweJlDSA1uDxFh5YXihWOfVvRMJb1f56jOb71osSBDL
BYx2gK71Cgh0ZmPTG56jAF7dhTDMY15aRXKcwrQdxlvWZw02BttwA/vcvni9JC5bwSvsa4TITWzU
6toG/BG02nmyqP2a+kE/388R6uS3/hfsGEmU8KHmOo0MnPS+Q/P4FG1Nj4GoKyw/cSYQ/Joub7Qu
nyaePvzRgNCKkbWVt1yNGIvurSrkz/904J1fUZm/9AWwTiOD/KbbkhQtopEDBrjctM8kMClj7TUP
V8TOHLltM8kG+ubsuXp8vJYpI5sIn6yXqgDNdCIdIzYJPxkI2r2w6zFyJzJ4/mpPcfw4NTe4iV0O
Ds9KCQ6CwvkM2IRhckTX3arjA4Dlfb4e6LkTQPg9a4IleSUfi9zVDau70Ap266D0lA55+MGolp/r
x8n7/mrAN1+nn4MHgQOVaWXrlgs5ZfnHEar3TmGZNlDNktNKH1TueRmSh2txhgg+7oQsTriJlOCT
gCpZHM4udQhWhS0HsM2Mu4wVYySnlaWns0+nHvlWpFssFC12op5l538skXi0RuF6QhKPzKdhE5GO
3T3xv019YGlGz9G56eQ/zdvABfZ0S+t8v54ZoAuiEmMoTZghKkHKZ7ldVx2jW8hJ8DQX7hhHfR3f
sXYVN8NSJm/JVvRg+0qDJoils9Zezg/iXsbEjyx7Qqejdpydq2gacL6zFyG/F6HDIs0LSv2wYXtF
ZKuAL33j6fSNtsyHeJ4TWk8r79N5X3VbMkIktEE1uuklquFq9L8uR6GXLmbvn7rI2C31sg1Fd7aS
LAdDU4XpuxzNaEMv1W3Q7DLHsOkveko/3HDxxpX8vH9iZmwKaP6szajWoVwQtUdt6UrPuma6K6Br
tUCiXasO6trHQK7//Wa2/2/7Y+IkVONu6rUB31zLk2N2p8FCHs5G8ljNXcPT07kRtxjq3fyWhikO
rDy2JXuS1liO5afsB2OnsMhIbs5joRQrNPMbH9jDsToT/Rrc88bXi1tqKb+NAEs0fUawVCpkPrq7
MqvmDJQAJw4oD7b3i6b8LMVFUzjgwUvWCbWi8TJyG92C2BU6YjTcYdux+zq8K0gOwo67dsV4iBQ3
vgRZ10fsSViygi69NX874tf+dppYKhDyiojuAu18U8/+3qzUpj7kHFTc7t/zI31lXe7Jd2MYv+o3
11Ddso7iP/0ClUtxlfJw62tKPIQC1rwE5gFehq8cbLCcpgevFkVSVHcm/1VpSvs5DSSOEbed1G6v
RFUny1Gi1/Ra0taOJcx57XdFZG5jKIA/PMUW0pvo+NPAjxjZxzVvRgIGQv0tTUa2KbWlX76wa9RE
hcrGuqONorkcnYa5OGmDCoMSiFfo8a1Gdn3s6UqIMcBKegkk3J4sSJjoEDA1/2gO6CYEoD+3WEqP
N3kxJwf6Uzqa195G9rBvrnjo3H5KUi4a48sjV5hD2VFjXfrOMnIBvTyC6TvRfP4F0iDg0SDuev99
S4Yow+r3wK/iqW/qGfttgYm6AfRawvEFsQ6VnCv9IApoEU2965Wijf7Q0EvNjasD8amsAe9sgB2v
9Kdn+FsZNizYfygWPrvBSB6mAA3X3omHN5XmhR+qXnDNPpAHhsg08fWLowmfE8SlV3yavDCwKYEo
Qle7IuY4q4oenofp7bqPYc4Uy+lasZ/ZRj+yeH8TH8dhFkkckBhtFLk3W48rCAVCGHC4VdAAiRM1
Hw4W5UmMTsRGtVauEEzs2pa15BidpyV1MTG0ythJE56/kzwfJko9xOlliTE+/MBxJCco64qhbWKC
MnjsCOyx/4b4BQe9XmZf+fR9XsxOxFzX25pEs4wHXiskNTnCcO95VyElbJM++3VUVv1OxtwjLbbk
KHP7G+KcA5gxxyUbZJiPOi7YorLHf4SxMwKCi0CCEzY00v8Vqu3b/FXKnvmtwwiZ9CQ5nBGd5XIH
o3/cg+M6y+bYAzQBgzD+wZ0uH6uPxMOeW13iWgaFceh7jbdgwaJ9/uKSwC2cINjjABd0aG6xy35P
TIv8QeEEtmBjirAslIeaoAcgHjYS/CfVwejwa6NnbX37SG2DdjZL9DR/BEW01/rwy9yvH+hZTMzx
pISr0/Jhu9zV2wk6rtLK9dpVRTgeRBKTEytFTvDq6ZxVpPvmFbt87L9Jf0vj4DpfXpWJQIYPm08p
qI8nYcPcmxlSX9SNUhuG+KfMku+t3MQEkSZIKZTyOHiP0s1iYfnHCVFsORzxhvUQvjaM1YD/rn1N
kzMPvyO5hvcLfz+KC4o0NH1gq7hEjJw+NGtmYktU5XKjZRBFyMWMTAFKAGJmSUH3a7ajIBW97Sr0
4cz2ZwTvCMDigq8ND6n39nXc23TVvDMrkjm9aYLPALFWADjzFO9LUBaXYBEfuoCBZmizKrmARE7Q
WxOmt/YkzdJT0UgtsuCk7wClc1Jk0fW9aFhEUrFlxpc03+BG2NZ6AuXoJc6RK7k2vXjLUqCarVw/
HM+c68/x3py2fT6XhsnYmHMyanNCDdKYMOQs+x2fLtSMIJ1is9HpCwZxVhrCErM4dPYWTL3b+b2t
In7hJkx8bku4mbVPUj/KebY9QHwqg3WBUPMlEBUpnodBr163kijo5edD+KpzUxDOpxxcWTBxFe6m
h0AyXY7JWWypkEQrya40lHLQFbDBo0TA/to8aK4WS+VOXgORC76cMy2WAptUE1NP3S9Sglp+9G8Y
81FxQjbxFprsbY2RY2abHGcyPMeFeoR5l7zjTetygdLXynIyafTdI6gl72njKbuKqjOziN9nbX4j
Nqy6yyqgDb7aJkDxgaYaeAkqC2wAqNHMeQqc5XWxquiTnkWKvhUaF/n0/V7sJ4D3nufzqaLKauGu
oetEtEL26ZUNvnz5KuiTvAapHHhmn7Mn1aP7W0ugEeV50v6d8KQCiDFFfTKdmri8Eo/MCoHRXlI8
MrGgAw1LN3AO/AlnjuUcJCYPyOvFpi9gK7fHzwGJnGSKkBBsafK9gTQwl87GcCN0+veut1ZkF7aW
u8PS5TsijwOOhtXjTH3mcqNTalK4aIiK5kE8OYosGdiStTc8J9QzsDbtmxHgh5BGykrjlLleTIrz
gEAkJovWCCP+eLEGQAEPhL2OSHLiPF2uUmzgvkWma5Jjci08K0BOj0kuBN6foXUgZzWLuHwzyeue
ZRZIvBwniupob0iw3BS2CYq3rgjInQ/6CDMTa1583ey7EGoZyN3IciSbnsZ1fNW7m58LzSDGPJzM
EOj6NPhmspOLqmBXUdFz6gf/UyuQNUD/AawOVb/cCQaarC6sVz9I57Ragqzm3Mtjkm59vROHwezY
D+5yldqaGEJHCdmPaveoxtf5T9wM7dtfss5c1FMSPZMwgDX4vSPSVCk6fgkE5WxFUozRq+7B+lEa
bF2CkJ82aAwI5ul77cWqO63A6JwhnrIIGsiQgOOaOXeCft6BSKEi35gtVpR7csB/jqEAt2dJ6BDy
OhlDvhRJJdBb4Cn/qRBzx2iSDxD5P9yVZr3cV2ifD//b2IBXgDHV7Uto1nZpcUYqQ9fAjHMhCdN5
rheAqqaMvePfhCISvS0MkUix+sRFdpej+aeEYLkWE2HkkgZzZqMARdEiTmykQL99IEpIB2Fq//mB
Bsoejo9l5vBHhlr4uaCyOEfcu2I8ZhNb6iAmRYEbd4+uKMIxoU/m6ALPm4Oz3vwfBPELIBUeC0dd
3egJwdrbTHg+lPKJzl7MP4j5O/HOa0qcJ8ewcel+hHPiEx1GK28RpesUudpmwswuGPlWbFk+bN+y
ScaV7onkua4ny575hJQgUK+l0zP/vorbgFcivyspHbPB9XdCV69O6ez2x9+JGMZfcEmQ2jYELapF
iKXmHjNDPJwJ+o49qCDL62v4XV82jx/NYIDKprR6bkFigqtb3LYDSPHBFkFA9REYLLn1o/4M/5+w
uo7Ax1yaji7xQRxKBU7nwRssFkc4WTB61u4oHmQTFnXNViWmN35OOq/Sa+Do/K2K+FoCTv4tQ9gK
vKoLjpuTfBqlTxthzSZOcBEqvjqFKPwbLJVc/FTkeTjhGaj8Oew7eu+4xtfNvrPrEbcx9zzvRFMJ
qSC59un2p19ldWrEf5ttMzum3rwldAdsMLbe9FLJ21P2DF4620jz7ARZQOWtWuxIWhY/4Kd33Whs
sJTkzWNIheE85FARQPtINOOcGVkcT5xv+M2HshLbGHhSmSG4lauFZ84gF1mq/EnzZDAg79PdaF5Q
+/YrhhHasu+BtVqQma0emXg6jkaIU5snFsgfhyCbedZ5j5gTCdjEvZENaiYesIPqiDYg4llXV9Fs
NcH7HlnWvMVpiJYUbURSmTuzkBaMjvdwFN5+nQ+E/6EjB9zF08x6UEJHq/A2X3bY72/ngklGsvef
AQ1fTQ9IRluwOE5qmo0OqZHZf1HM/Zy3y3JaTvWK1IiOVg4i4/rD8ceeaHIrM/KAQKXRjQzFv2Um
ThDTFdul1nl6oPyvdV31tN9M48/rPAMx1QFOhmajh0dt12hts/WO2omX+dYUgAD3++uNZ3R6AKOg
BqWlRrr/w/MNtRqqypWyUK/VgkORFCHUmwp+lbZ6+QExUc2+jgNBQRoEuWUEIiNeJdiOCrR8MuiL
0qIP738aksSLRqmpKgV/PrYYJtWWShyKMfatu02+bprEROxqDqYWhHklO9fS9jlEj+wfI9wfShMR
Genv3cSGFTpzjRPDTisvLczkylauOvmyloHWDfmu8iNwAQ481KCq7Bx9Jr6xdq9xwfQQON+bbBvN
GGJk11UNyHp4XU52/kK7vqrBfX3b68EuPIS63/jKP/0Oehvtj9ORIq3TJcw7QM6kBXTwSXqNHnn/
onpwXibIWuOFEq+eRmns2CgTslGFNEhX7T6seKsogn5qDYcZk4psa1czvZU+RQtV2KmlnfdQkDRA
SrxMDwwFe2slP/aHR2Ha/Rg+uoSyzvjNKhw05ZKLPHdFeiYyqpEAU4/07oNenjur8BItifQW3liE
bmtv+ZjydJpJp2P5+ZZRPJByZQdOJzvpw91QswA62H1KH0FRVfCHS6tObTOkWvBTzohnNAgWj6nY
q9yiqaZc0N/HBoBxTBrFmzne+y6aZiryeKkLg+jMOGThPkuayMp5lgyUM/+mTZYpbrach5VuZ/yz
wunomY98Ln+46X4Uqz94+ihEiGoFoFVfeG9HNi4hb47Zak8cNT4NVhuYyBvmzqJUrZazDEB+JTlv
z27qlGBR5YpKVOzYX0qq3g64ArcPqTk7jSWK1W8zJObqV+/emUaPLWVDVlD2Z0vkHrO6WdFz4L1v
u20KqLYs+Slr06kEhlrxPOVPmy8zErtzxaJbMWaUNbZB4B68sTzAlyDIQdY+jTVRlzXWo/+/0HEH
ScrAe41nIz0ex8ltcd/11HsZfavZCqrog8ljrji6cDDPz/9yshfohO6mrw4TMFoxXj+at/hFPayK
LBmjDxZ6u0coBeV+VQDhQyEPTvNXID9xfD/PHGMHDIby99RkXt1+BVjDAwZQL9fsBlOn3qltm8nA
uvDsW7aBGPNdiyTeKmyh4sBP8QWT3ZDT89kmmQRNm7SaaXDBg/CXdC+IPPsoVTVOQR1wCTvuUoYX
KiIVegEyk3PNH2DFSsknQO7LS6+A0PU3ibEvK1q5aU4twtcXbw4jv96o9d7uyhuwvyanqhmR2HTe
lqGC4rMiHBENM0LuJRk2JSA4iYirsb/J/1NkDb0xaU28Eadi74YmMzm0oGTVydl7c4JL1MkiLBk/
N7uJ9+ZNHmPJikNmWSLgi5ocmbplXe9iIoeQaFjt+AKNOr6hFjQVxuSLVrnnbkam33LyjC0DYCt5
XTz+5hlFezagp3oTZlAPYIy7RobZl7MpBkIKIDwDKPcvGllVSsoPDKx5eMfGT1pK0w0QplBfohdW
7s5FNdx2Z4GtK8tNGjFREvJkPfqjUC8Y9fuJ9q6/34Qei1J73m1B4Uo96d7qZNzRS8YFLXe5UQNr
zLVQDAlvJJ8TvG8+xLuQck9MoBSpn+FKNyzxLXwaSC9KbcjUKS312PXhb7m9N5LbDSCSu3NvPjT9
xnKEKbXhNLzBBTR9kXtcyF8kkLokZeIbYtrm2co8y3gwQqUOfnW5D5sIjiAHqa01aYGxbLqejO7O
aZEboo1YI48XE6EYk5I1DqMFYjQq4uIvi85w6kfgWq+HG4zQBquy8dyZlKOG1s/5YWhKExllPFrk
wqqWChPoDZt6WJ8j2lj4OXZcgODiyv3zbZcmhvNwmz7UrFckO9osiDjS/BvqJZhQcZpFqdFy2Lo1
MRrAGgvoVRorAKrNtaNkMSlEIhyduN+sxHBHq4le21brlmX4OksEwTuNheE73KvZloBtwdrByfFX
LIV+FtnCyXAM4WcZVx2hr7w0qZOOIGDJfJEUxfW9c7FBteUXl983BQAioNHKtSszX/Y6U20Av85n
lAd4ePTQTbRmrRS6If0lR/bUm0gfuEVf3SIEO9wXMbk6IhQdfdbKJZHrkq1LLItAmqOm5FAfhyRq
rA1UGIv9eaJco3FrkUQeGy152CmJ1m2kUNAuuLlN3UW8pDx+T+r/2jdvpJ4PwhXF8sZAuIWnJwlo
HU9shxVqheFFRc6QWqR15jtkA4on9+TUWGQPkTbPAjl9Q9VKulpikwKIB0sZ1qcPlJWM8xRFyFBv
pdeIU7ZdNGAOYnNSNJ1eCXRbFbin3Z0C8EAqhIFSuqQztUiPc7Be7DpJx563ghvqEvbK83aBRPb8
aazGLPXlisGCjgS7RghLu+wH/VynWEfd/xSWUzfjm3tqhGLN+ums8Mk2qCs8/ie9q+cUZPSIIx81
RBQpmX69wjYja/v/JexQRALdUYiPEwB2i7Uh7uUtVpbeMj5RLMVjv1vgucuoedgL+/hapVjEPp/W
0ZdJ4O8KAM3c67owcNvDNBZ92jn2drLAaP6H8lkAHiw1KTHl5IuhsFF5Pe+8/HCy2Qpiwqp0rjwz
XY8EkOb8uiUBCKu+pYqUvt5JU/S7MUBKDI6kUM1LaiaqlvF7+/y2BJumB/dqnetQWo6/xuEEqyJB
5nWtFl04PZ7ZzuzE7hpyK3ipmpDcT5vdojVbTZJ9H5yHekzlFbgiUgHi2uAd45lKSCsycv4F1a7y
RneXrjMNndR90vUjQ6KCX0yJFvXly6YVU4kAb1S1wfjOJ4+SXcgJLtCkH/a6zmwZYFF05vM2cQ1C
RHUB9/dp/DEMz36lzd1mvYMzHOOhGMbWiEIEBaYUoGQg3SnWAvckTL1Mjkiynq4KzLrMncqKvvTy
050G7NlOOUjqcGzD9IBfdtrF1vXw+S+3KWVjAy8sKar2sQg6C2SGQHvkEkXPB8hBopc+nhPB5k8n
dTL/tW+zodwnClMc2bXqu2lFGU6Ui5hYjwLjTGDwsYacbtJ2PKu6CctlpPsea34Zy62LCgKc55hI
ZMFln/Y4rdHYQ7RYE7BJxMW7HfVPf+SUSZ1iOxJCgM13hzSl2S39p2hhANzP62iDUV1aBsiyvHUn
4lE1YCMxdDjfqw2yQkphvGTCpo9BCVV5/4VrwfZ/BZ3yZLP6gMnzzGNCFJzLJnZl2NwZWlCuywFm
lIP/mu0uQPPYa/PZ2vAHdmALaIqYUfTBo468U/KhIPlYX/ScpPne7l+L/8Z3XpUx3DOvX+D9fd4v
3Rlj3ONjSpRN4oxU+I2PCeg1aDD+/+lh5Ht3amJ1tgG8sXwLfS8SG4iuT/07q0zFRrJ22WH+Kepi
GeFEoiLGGSMC//DD2MLF6ju2hhWstTrhV1VzvZSY7fFXnSmcz1se6Xm7B6Pocem0A2RDY7opUpA/
OY2vS/oz6pH89IEikCsMBO7jjBp/td8opCmUI38RTl9MZyw+4+d9x8Xw/LL1v5YUVmjBZmo1u1sZ
LvLEaWTU3wbMLa94WPAdgQJJUHsdedeH+9rfpJt27grpfuOEnGF7OA0k5PkTOO8ff7zU2IUyLGVq
9viOPEbeufro7qzj3BF9K5k4trvbATOh7/1Iexq+wAtHjBG2aMbczn/qldsYnOql+Pldpt1Dw9n8
F0lJxQNkPrzeUX6lxKnfAoD7ax+kx4/RBD/3F+s/8s26qvG5G0DQ7/tR/V4aQw+pzkfkUv66cLNO
kmYwQ24TEa6x8ttQ+EVDmIH+Y5boWD2RzAfc2KX93tHxqJhxbcM/SAsdqJbdo21YegQ9+ZSQVMb6
u7dnDDx2zYcCR5rfQQLJK0rIDEwmw5Dh4EB20qVcgjxn0R1lWbl2VP0HP8WLQTLW84i+XjQMHQgX
vLyekQUeUW8FCZpCX02aEAi/N9nKtOBTR3B9HIOGQPiERgOM+cqHRVUg13qePOSxgbpHuY8/kG2X
ipZ8LEpGWn8U5Q3hhYQ7xClzpeHKbHuZqNOgqesDpeoyF3kJPVqW4pi4f5S9EZTzllNxft1aINKl
CzM0HiC01cGu3wQ5WWBOew3cunfcVFU0iH49MebHLkNwd7OTAIKZXpmolf2Yk9DLpneodBhyKtEN
FhHo92vGLS/IxcSZT5ikNTDwvQTNXDZn5jefdn8LhSMTTz34veOL+H6UzPn3kNNr6eE3gSp3VmeV
oNi4ZsWoPmp1IGmDjiJ+cECc0k+fTKqpFyX+Fusnb22DpOtoyS+2A/Lv8Bo01v29UWGcV3bW7iib
2SL6wl0R8IWM3RXXf2E+Mp4D4ZRajm6cWpCGXetO4j09RM4bmGA4RHe1UiB7zc2lYAXXirBXD6kZ
CoORqbABTGGP2ODWiKeKPNOoo8PK2U/VqYHv1DIax5Z8tdhYNJIzK89dYjhc0t7GjDvk/nDET7lF
JpW1xtvsEHBh+rQSm+GJQ0xCPye5REL1YBCn6a0PovKnZVkCpDsbS5H+j1NYDOSgv2xqYvWv0fJw
+oPRP0jO4jPXY6i5BnszM/kCkSE2ECJOpUMkNok+PF6qvtX/YNo0BmvcyOdbpN0pOtqWmi3xvPBY
xv0e0ebGdCckXgAnzQzVm6a01rcyNjcf3X2mxNhlogjc0emqGpOli9avqwF4P7d07b5gHYCMJ6SV
6YcJ3JenuAja+8b7DpRNldqU85pwuzKS4Tkhj3o/Awuq+dsV2s/iW3xYMwbDF+jEKWMDjBpc3WRz
KHhxBvKNQLBMjydRmYiIV83nD4bw3Mt+ZQICJ/lNsCabRunZom4qJtjZhd1p19dpWnJ6iWfdP5xn
v+s6O2LWr80jZnISHll1/s9s7rG3DE45RU7s3woYZp09KsQ5REi+6Xs1EJkHot7NdPM6kOdV92go
Min0K3kw5559vV5vbq2ZyrBGQaaUFqRJB/jOTZ4jWq/5zoEh84lZooqUSA8ucyoP8ReJ6vhCK4FD
pwiSg/ChWRz7t6SNmOI1IddhnSHXwzvDE+nyHSzoyfJtJSc5/GRQfYLiK2TahuSSBnUtChVRiguG
7KjE11saODTXCEEXtj26QlpWP/pD6DxLJgJwulTpbUzt+u7dvXEBLciVNB+wOyTkTt+PjhSh/t99
6u+hSteb3HY+sklvW/oZFxtIeVf2nufD05LxLQ5UV8tS0ON0PrBm2u58gsd+wGW5Ny7w8gx2BSRK
zi7mYzK2WQ56s3ELR17qP/opvybB3DWcgWdoNk2GQIlhT2FvKQ9+KVnmza6yIjkNRpEWSdzVrJDY
doYJgW+nvGrMorje2m1r19dZGaVviXzy0LaycFnRDyqr93jWECHHdKOxbcVebObpd8bL6V2NmB23
tXXriXAfw8uhy/WsFFRcEFRSBqFB7JPpdeJexNCM/33rryQ9SV53WZPqBanjxDyKgtPMexVhvxc5
4rs3V/mh3M1gHwzWthNswTOFxENRzj8Wr/fxlN805jm7y3sqcDVeQUC9KrqWkBCWx8J69SXFFS79
9HvV+jT9DHaqiScma5vTAQ50VnN/lFMeAjO9b+bGKDnCYl+kU8HgDDPlQC3k/2my/ZS0r5oIs5sE
BXvpa79nxRPFGj8NdYHh4hK56ke5yvi9r6ckHTbxE/BEdXOSclazpkzKCbjbZAYUc0O5Qo8BweMm
r89f5hH6l07aYXPD/KNpK4uJ2tjiiTa/v2Ad7QJ42HBgdUQZhYVuxjC6USmi1uDQzW+UfwaIhipQ
M7GTcwU5ncNhrkfJFe38+ponZ1aoy2yd3NZK0tWD2aGyTFI5kGOpTMyXuYH6xPvnp0SUMxHQ9o9B
MV316Zz8pQduh+A91tidgP33lnu6IklGkAQ4xXBtTUDjlyj+f90I/SlBskidO/blIsXNe9dIF8vA
bc7QsWUIaHW3eMJN3b2+DYOoNnU9AR0dxRjGEC9pqzV+YZXcezeu6fzu333TZh2/GmQnNBolOpd5
uda/YU2KWyNDvGCPtL23J55p+P9dP7QtekSU15lpeGlrcO18bv0L8mDEtjIGIWaNcop71otdp9x2
zx4FsCaIfBd0KDX5LimyrP/q8s0Et5K/tJRz0BQSvG/dWEvUZBeiHkhCeAxd+cxqWMfDEtQiSKYa
pH202XUKmMfyt86q7twEINseAmFHr8wOBLuWR/t+a2rTVknZJ1rrbdbol3RSC5uvUlVM/FqR3ovA
ojvczFqPB6rrFtrlEdhlpqvX1lb6mkiGEuJZERR9W/5dQKJHwIB6QCLVyYf+HoBqLqhkzEj9We1y
epovTOEEgQA27L7AqqcsREU06v+G9AbKXVvlTtt2YV3nVBkru0bo9Lr5pIL8iTJ0OVBh2wCxxft6
0n8UTinJAItazPm+sF2DWP4DaV251wQ7cpEsO0UWMy1EVzdGx3zvF7Dfn/NBnN9WMHLDIAPc9bWq
xXzdPqRFn4P3KJYu8djTa1aaJDrVH8GQmHE8Ga+yCoqHViUWiosWC8+wW1hXCxoUd9IhQlbWdl+I
LLuMbOCn79+M3EnbLMkqvNqUSILykIs8F4Jj0Qb3KqkJNP60LDo74eWPYwdcQ0Nt3M1T6hl87ILV
hW2rgbbDQg7Hw1EZh0lFSLMStR6Ufx2g40Z1rzBvt247NOVrTYdBTL5yTzTMVQi+zMYcX16AYwkD
sKrcoFZopN+fgjvts/2a//u8YBW5ZlMXYk467w15HIhrdCswmXflwbAHVEhJw0hjyo2s3BhEAch3
+zHgdCw4/Eil6YmNyPu1D82GP8mpk3ORKMAqO6kV4Vrv7/p6PgdhEACWNAxSWpX2YCRZIu1LGYYn
H93lT27gj4Ci72VuODxGaBewJrT4+Zk0WEnUHsmGV4eM+twWYpKC7G6CNbDApoxZ9W25KcHihS2K
AUELvj6Fe9R2pGApJoc4UCWrTOpQsC9YK7IKyD7iwjC+aUdDUGod+94TYtVb+Y3DarElp+J/VCbC
+xNAmHYbtSBm6UXza1rFbslopihoeNupuzojnXzB2GKLNMxCvIy+6jlfutnp3gG+X8ckOJ9CB+wi
cUxV5Vr+y6ZHY+pSiYcj5tkD1SUUtG20Ju3NCwPTPV1yDNGKPTXty6Wt+IlS2sRLn4NNdKipHIzm
ez9cEShmo+kEdG2VrInppuFCl+6/sssSf6ylTbYjcQ57td9dq3DtgEHXk+Ha5JrB6kOsgJdwPwwE
ruFtW3aFto327Ct+S/3DmrHEvl8TJsC54mRKrw0pcRs2eHJvYPC9H5tXfxF+AcJopUzeqQ+02OZw
5iL21omkcEcy8wp+xLnusDGHgpOFExo3rVg8QxbDl6qPsPkov7bRBPIZ35qcbXtJ52h/eTrysGB5
dKQyNJ6fSN0u/IFs+Pzk1tAFVO4eRp/q8V3pg3qWGTyCqo8iYEjI4XrbKy7xM8DJW56fKZUj7fCR
wLUhzGg9JRHXNv++eDjvbQ/CXJxyjGu8kdjdl3eyfpPumGB4KQSTn0p9L4W9S1rQzJSxh0MjqTE5
mEMAh2SatAC9bP5bOFqrf87Qrq3hzUF1tdvNyXvyk1Cc9U0TMA0D8aTqS+HuIy6eFE+yl7xiUDGb
5lzJEXnh11fRfFalue+itDxAlKU3RkAtwTdA+RbRMePlLLAytSmaMw5+rLG46dYPTW9nVn7ST/eN
BEWoFmVNcO3/duJNwPni35pljPGUfCRNQzNNuj1H+GY+IpZIzzWBNg2XxZ4YWEuLJqlVZVnlYipP
XrENPcN/qFDO1VM5gZ6+TcS/VgOaDfw7VllgZJRqSRKRd6cx1AgMBf2fd77eLgUXGnHGNqOWXKu2
oJSWaHENESH7FdQuvb/0yITd4+iQ0Em4JGqGQgCADeEKQxDoDG/gp2WjV1U+TU154AWJCiRCcQyb
hP8+p2AUeMdcYomL2g8MudnF2lrbDxmUJWwKX6i2Bqg1qI3IueOMOYefyerFP22mJk7cQ24sfBwS
S94eu9Zsi+A3VZd/MfovLz3jp2BJNU8qk7lj97cRWhm3KVFq0rKYNFRQTio7drqdytZoeLVrDiBj
hiunr7JHzJHTWQtycQemG9gCRJGYmzU8bJvCUGZ1H/ZV2oISLczdXjWOxyP0UUkg15+0C2oPisdj
yMlHRuZZe6Ouv61Xymm3JICcANfyEoi8DT8V6WlJh0dDSQ9FhD/pVRENwH4zpv77jCDMwqkb+JAG
WWm/8cLqREW4ukQCAoIfvnPgCFe1NLLwn2KjH4bnrax6NzEpOlBCHfKqn3QfZ8dboBXIclj1SY5l
OEE7flRn3vpbXb7UHNEJ4MpJ9oYpCZOZbrU1LsmEV2H7a4DgfAc1+OKY+b4csKLIXRI/JD+jfOfx
hmxziTpzkFPnKhXUL4ki0JOLqfWJx3w7v+2cnBgkag4Cms9ugw9FBRdp7ye33kkPj6jjRCEx1v44
h1sQQfqGpjr+y57VsEXwm7AWiAHuac/2+H7VALKLHWBthJrhP/0NYPttIE4b/X6Q/adGht/E4imO
Ik53x+7Ntxh42dkiYPqPBXKCMHS8SZwm9NuiH+rnP3ealkUuy3rq5B8B1MZ1R1FT2a02IR/6owjF
9t934FJr2uATyf3cRn5B9n444M1Y6IXVmIMHB4DlF9gskNOvonx6kWdmn50jselbuDoruGkhgOJC
56CgRrLtn8k+//FyB/GAhD77rilvz9qZv1vl7AEFq62SCSyBYq9LL0e1RgQpXxHnNIhDwqDY64ih
5ZPKU4KA/7u5EU4lyTf9CT0Qgd8qT3FIQFKhxdGni3JqN8WW0awJtgNRkPyklL3Pk5VIfPhWBvbS
uVCWeqRZeOP4+WRQpbbU9lAvKNaYxbQRQ+f4CrWoHBDxfrXtGmpvoMQRgh/LPB4sILto9FDG/kYk
vtP7vCX2T+8h6NdkZRg6Iox/7mAEh3ahFCwW7ru4p0Igarsb83FBU2TJE/9GnRWEg/uokgCrJDtu
rnbEamNuysz7VhXjEdiPQUdvcfBFFXM2c34HEW07AVFDZHaeoCUPdSSSaLpk1RAmkaormd66g0xz
g5Dgu4kje0IMpUcC9w3txrAtByKcrdvSHqPNSWlpZB9VLCvSORxtYrk9ACstIBMTYx4BUu+mNsF/
/oBzKnv6DaQpMBjBZU7WkLg66fH3NpBLgHc6ObH6xjrFJiYyVhn4jQmwNchvB9dA6rXIrRRRGqUe
NhOkbi4w/zcwlPBTqwW/Tta48zOBEVCfCfTi5ULDEnSfuVQOr1sUt+wt/8lJNaiCm3iny3b2Lbz0
63yP2TP27DVD4XaQjRqLRtq1wxvR8Q7KuyZDCtJEFbWUKEHF381a2nfNmKXLRI4YBVVhKMsPBA44
Rp74wCP8jUL5E+G+/5NvXriC+oJo4Ie0SxkfGL3JJYiacIs4hfeI2fMgS2a+De1ptYtPTF1aUXLW
/HNAGlImglyRPAC89ZK7zioI7WDvtNdkQDgYcVwo5iyrzEsNqpADlev0vhVn+JTbF23wm23Iu6hg
W5Ha4R6Zj3DYySArFZ0w6G6LDGDHzhFBsDiwGuaMWKneuXg3gPRrtD+1WeSaVXiN7oPUrZsNlNzr
g0CRO/xPM3V/1zdRgpb2Y/4tajSlzPTbuMzYDd/2sk3EIjWGkQvF86NzOaYsryUa3ciezCEmlYwM
AiKfiRh8fJ4zmdNmODHAGdavKfzarFsl0LOFzGHtq9s/3KYH3RdZ8TdWp48i2oj5esNn9MgqryDn
ws7598okKM/qaTPY1sqyitLGhh5w8tPCwYcWRawJUrK6CCZTHVHMuEHJjlXudISGGQ0Wj1zIcpIA
PSkgg3dD4Sg9bSptgTX3rtr7Dr13CHlx6B3F2FHEo0ehWOEVcYOdH+e3xEPDW6RXENPSabJHcsK2
z/IotFT3xq6WemGeGUcUgxHD1EeqfI8g50abh6Iv8wfT+Tk5n83kFuIIFR6DA4/3Ob89cARGdTi7
uDIpZsiTgdkGFVs1bTy6SyQ10uk9AAUX/ndaP4gQzHtSVAMFsLAgRQ+6quKPnoEenoLVbgnZcxW/
Did+xTcjQt0uG2cut4gFrIRC1gMeMPgPq1aWIz+WNgtqJ+X1D+pYRPrMWXRtrayCUUy47x/CcZqy
FfE6TR4yDuMir9npIbISlsMHdAaXEu6CXWsjZ4np4iAvae2CU4UqZCRzNHPxINANVwNasCXzdHXB
TsYy2yLHQ7L2ROQS2KqsgwcI0yp6nEt4cxy87eyVEeF6onJk9k/HvMBuvrriEXcQkswrwLvI4+Ps
155j/jkpShki+m8vPjThpsGwBEoTQg6nr8F27+Oy2BH3lkwP9KdfOGT+D+d5/8AqWkAL7MzHb6PL
eHVWEAgcfqn4fbTSXd8iMiCvC4ZybTAZ9WWZ2SPP8F4K7Eh08Ctzs5SZXBN2PZCPtmm+IjsRuYrl
80txeasozWersykVQrGRSG5b3coYdHdYdhSAO6TxFA13ghxljH5OuV0jgEnJL2+FrwYdyYFrv3iy
xX46zZbSuegYpkNCEEc0nevVCx0pxvGmT8FBgoc2qN1mlV5j/L2M5+68YeGTaWv7T1DqNd/sZc7j
gmw5xInPrps5oFtTy/Xs0Jh8DLV6DbUlpLoJnOHxvzvTL7AqNeDQMm8FBZhf3+mfge0FO/93jJWk
zlfIgkO6558Q15XZFPfFGKoCpvs0bX3h2hYVcTxomsAWUX16asfe9632Neleg2AhW0iE797KpR4Y
orCR3SrkMC9neknYffYfLzpinO0FyskUvJ1NyfElmi4xWkKamgWGQuAJardNfcm7E7kicXD/pKDe
Spjvp33fMiBAWyFszQmZ7Ojsc5R0b2YlWb5J9P2oy6AwwFZMD9fOMxneXXTW7ZB+oWl0SeVr7Ycg
JVLg5rm5a00SxizPxo5eR3K7YnA3h0KJrxIeBJNELCokPVyPMVZ1g8fr4AnOpd7CKL6P4PlDlbFC
eAdOvfpebvV6QNok1rcnc2engnIJOjipKZYTzF+VR8ra9QKEuksfEAwSl8w34SXjK8w9cpiGK36a
jT5efetaYN067FNpwDbz5yoBY4fP/vjiZdiWklJBkTU8kFOVsjHOMd7lDkIhdLaElFvUz9b+4C9A
6b0EzuLCfAvsdSH02aO/S46flpZjrt9gEEXnOBOhrQfZT0SH9E0QOA5wEIpQviw892S/F1hZt7Hw
axostsZ7eblWcjmkMJw00sIiR3juZC8FU90MffGc9l9vc64FEHuk3OE0TD5kvHE1QPmX97eEMS5J
ZWzStP55DAJ3KQAfFQnuv2INtIIJHVSddPR9uHTCsKT8tmZX28r0vA2AuFzJVtcSj3evEwchzoC9
ZcMQ4DUPFm1YMWAxZq+uypAZcZRfx8qzKZ5r1x7VWn842unxd+nlsuFXCZvr7wNRwRB98fJY4MWd
CHPHHjUDGT+t7xpGRw7qrKXXxk6mA5aInT3Hbs42VuzFIlUSkDVIdDoCr37RDSXRLoMIrnImLS06
6HhTJa85FK/Y9h+mCD1izz8zz8YtQaRQNu3az7vlkyql5QEMwhJrBcRJFthS9SZC6ZKTeICH4Fo3
84fMQlbsl3YjSf2Z1w7QziG7Qg2cE/KFQiwcGdHUb29+/bZdQEmC+dVAjVyNawVDOJrRNVMmiUKN
cSGNWeRCD+uCRQH4pE7W8QEQHWr88XAAQ8HPHmZGgMGEggq1QxE8ZUp+um1LBXw7pppywzdQjQKA
AoMnt2xNUhH9pqWRRhbX1i3daS/hZWMzgunwOywmFOq8a3p3uikNaeiG21rP/KQOFjg7Wmxfrg3g
VTE+AZdOZ9hZNcqNtRi9jkvDR3Wr+4g9D/8POax1H++ORlVwaZPAoWUPJ6XJaQ2QdlkLE6Yt08Qp
YmjIQQqH6oBaX5TPic9fFI2OI3FUPWdeuMPRbi2T5mPwdNrJ3D3JezkUN4mj4ZSa3Uvk98lZd7si
/wOnzm6/w04Bo1TjWPYIVlPbK2Mc8QFTl4qTyYUhyfWLYgpiOhOWGDqO9l4TaMhMfS/1jUZp44H4
4X2063QaYPwwD6s/vnIgY6jbzle9nZmhlepUOhhCOnQ1yQuimWWP0W1gl0kTUsMkzcf3dqjeZYMY
zmmRjRsBG1S9QeNuDYnh0JR7te4jEEzbayliXfdJ4VxOoV4fOVrlxPB+PYcWHymeEUo13vnrxUxG
9aP606EH1iH351uzCw0+5fIX1950+O+vJ9j/LG+LwbeTR589WbB3Az3/UpHg2Cl6OcdOtJw48dWO
/LXt4wJuQskF5c4B31/MHPa8Rk3Tga5ou6xPcYnMOLXjFrUscX9NGOLUkxmXTb2n9b11NbL/lMwe
DVF3IhZtqaxw3QqiGb1T6DYsN/MaulpjXZvGCQq4FikuJEGLf5IV36tU+rKOaHK53zQS4qGJ/r/q
GqlU8+NVvVGBRhdIyLNWqaMreXn8LauG47WgzPMTao4RO7Z41bNAAyApuLVr8R9eV3Lq5LzhlVrw
jMWMRopbNZ85SOMpVpIY67J/qVB09pOXsbTb/lTKuS+1DH+qnkzQYrLni82U8NwXysnHYayiEyw0
MGI8HJy9QFIR07lEy0mqf5g5bq55++dT9swC1OC9AX6qjhqOBb3y3T1Rd6tp0NJ/xubvGKLMez3G
trtqu5oxEAB2bNprnE4qfQtq5VJtrNQVpswRymPn1xq4mspxaqYQdthS2FY25hgtaFJIrQj8Gjzv
9pfCrYkNmJY9RssQ35Kx/Mw9+H8vf9vHm5lULg/j/3/bzkouAUJgAx2msPe7ec0sRgRfTe/voMc5
dvbCqk5UiOSKWNgOTg3Ox4oN2zsqqKTHLV6grgmiu9IIskceZqyYp7t34sWh/6CVNeRqxGG0mONS
f/g3TnWb14DbDj7+hVAJzCGKgtVrlwgZNDlGV4C85K2t6KdZ+SdW5nfYMXsKiGAKU/KCViX/jzH7
6Crglf4eei9vBlD/8wnQZDFsuoRvM0fruFYFS8vJsm/mj96az3XC1KX2brvPifqm4j6bBnARNS4t
8lseTeOtgSREvQWRQTg23Zzu3NcGGgMmUT9DdE8fDeTabg2y+z6xbe/VeooW+ixFGMwAXRCulGZE
e2HSPQFKBpPG208n13GrYLa9odLXxhyLvTWhU4OdnpWc19o5P4xKuNhyoyfQjPKMUOPD8Cwj/MRv
LfUL/UhQpqFpjoxtCDIlzMPXLVh8Z3I2XSFujVRm+R7Ttnwa1Mpk65YyXGdyWV/mY+e3NzZT/b8X
ekQOCHd3ZG/1+9WHVqOwhNqzhjH7v/4bvUnOIgg6HANYZ0EeyoOlEFtiweGDLeOb8Xq5rhVbvlEi
EkParQT/G7zDSZvRcfgRgR5YwHqpXG7QhaCuADsFQ1VM2FL4tH2uyAF6AsUA9DcrO3KMP4ad9Oa5
eEAj60ACVJ1WqjsdOM5wbbMHyEMmiFoIhqNARzbRrZaAhTVoBRhD5Ag188vad4ZxbRpoKs3z48NY
eK0Tc3HECCs44Sms22PfL3jDP9w7ZSt7AfPXE9m0I4MYfVJPOGk2vvSMRs8yJ+CRbXX5PaznHGx7
6GSy8S8NbM8zSCPDdoHl34FWIf2UZFhn1wNcrfrQZ4uo9OvBQ0DW7N1chTNCU24cZzid39ZjgG44
ZTQ1lEkmPvRZS8w41fo33ob+9qDEkqLOKbM/VerxlzM1DT7/AqD3LDGidVVL8/fpU/mSgB5KT6NB
MgcyrRBvrbbvILV74xucwg8HvGd4bsxl/fwvEIfF+SYflscBQp3BDbrJUga2zEpqphEWJADZqTsq
dO9h2soWOJ2/mA0aTqaeFE0Pr0lWqiaXWCNLW0P6zCH29ZrjlDIdlzFnFAIevzSaTsI3tT1CEpzj
ZIFbtd/PH267/4KKAOaualCwPXbJs9oMfMbj64ca1plRD+ajSnGYTK+uCaPf7nufEBSXcx6blOu3
LWNuBiOMiTOWgZ5gXLOSN0l4zMtYOj4rZZf8O9kM3NfKDjpnr99kRRgNFnBGL8L74Zn8JTQxkBF6
rcOKNtFKu5oJt1BsTYrnL0SlSXyYjee/2nBe0zruqi73PTVZHV+LXyMGCu+OrOSzM3bGZvAMYQ1q
juOW3FC+Ke8ouLMku3ljIfbz+5u7Z/y+4PJTjAXjqjySblY/fwTjtrfnPq5GVRMHYGFn3d8omTvm
W4zijtv8G9oiluoOZiIOOwuBtIODNnv50wF0OmJHJQkAC0jzLz+ZQnaB3S5Fpuj7NdUkIQvnvFkd
YFiuTeBamRngLgnCHF1JyAqoSom9UA2zACYm9xZq9MoPj/9Amk8fsPxeEf9y6bR6YorF62Oj1SXi
A74eOFkntP7DzcbV854Em9b5ie62t5U1t/lGOPiYYMygjZsyUdosj8SnCUx1CpfC0BCJZTIgNsTm
eUe0VfqycEzz8Vm6vm3cc59T+Ohsgse+WuaZWuy2d0LojDXwvO44FP4WA2OCpWb5nASkizXIXDt0
SwuXOM/ECiWPTdtsy4hUQKKlFaz2FAhdxuZRk5AkjRbbR2nGsED+VPU5Qa4L+U8OaRjyuBHYFraS
Z65OE3x4RaEgI4JbVWu72IvRpBTaaaCj//6TDvKppg3RKHMv40amMnOTSiGJYIB3/JpOY8voO/pq
vxK5de8pecdA8JfERiKETqXhl8RBst9nr3j4Wruwc0ncWGJgmKJoSUBWlPQxeoV1LPaWaYOYYBjj
csx7NWQCDS2a/j9Qy+a6482B8xs9BagDprTjttIpqxeur/qNbjjIdh51SubVbrAhPjFtvoS+j5+v
Buj4W0rIfHHOc6uWo32pd2hBc2IzP9C+uG8u/nYAak9ZAZwOrnj2p8eH97fRcZUN6eNLllvLxcua
iCNBnd3NMCBaiWDKot+w/FkBwyitlm7Ja9QR8lC4R/eVGtFD61xCNxajfDWBQHOHNlFHPbAn8+5L
tWLy+7wn3SgtNFWzDdRJPxtQNYY4Q86nmwrm0+7lyr4ATgU9+Na3kH6nyLP4CvV9uByCSQHXEypW
pTows3tHn0NHOXd4LONoOhyCnkJmC3ukAT4mj753ueUE+Qr+KEpT7wppIAEUwFPsVFjIyep2XTjC
Vkx+m3nzOCITep6xAw/fQc1DEtg/CLn6YMB7uSEHzs1FnRul4fl6duOMcQ+TAtJC+VcO8HUO4mMO
KuAfvpD7x+reYF4fptc/SvUSuMlS6KQ1Suc8N9nkFYAVl5i9g+dMFoU4L0YEP9QaFWXPxHB1+bAq
yMRTdV15aoP9fbcwHTgS6ZWXReITSGcgDR4JNKa4tuDgbIp16UbmD3K6JDDdi8QO2n771DawBRab
l6nbvFPui3Pn1QbCOJTkFs4fJXpVtiV8w7u7M9eb9lGuMmoPEVidmVDFNHPg6Gh02UIwMtA5ltVN
3dHiGYiUHe9pWNvfNV+vxShCx/aAnS8Poiy5AcDUzAVMIRs/ivTEpVejS+H4iobnmFXoyPWtDSbK
YgUmpBD0W4Q09j3hiFip9uQRw94/bFBNgcoqFC29dvodNm7/srdEbUx3KgKPa0yzEzCG1Jdww23P
4UHgWNk1UuUCoFrDBDjo+9xBDAw2LQuXukunj0tB5T+gPjP5p/03R27zUprUPt16seM=
`protect end_protected
