`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ms6qqppAk4/HrFCTQ5ZNL+e3VvC4XPed2w5Hhua7yvyqP1sb188c0XyU8La/74J/WjBGJtO0wJwN
kcluHuxFZg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IfD22Q4PkIixfguiLqLQwfGuS533W0vLscqGOgLQguXKJ22uAkBjuCyu6ghazvg0kS4mfZocs4rZ
inkbv5dEjPEPASsDJCIZwLTFua2gLTUNOe15MKHaNrIdr/t6hNASx/u0O9SyMhLO3fpFM4oaAsCV
GAZp5m5HAnjF/d5wAys=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XPzqNlPuJhFElyAL1Bmyo6okmNwej+KGb/8UcGD3GvmAx6kk3X8YeGCgePsS8GLaH5EXy3pEZXj6
5KrxmpErE6HlUXVbutEDVl9cQXkkD/21lFWYrhs/RMEiuyJP3dNVI8ET92RcGjgOZTRDC8xIpdtg
nAoefFsZi6q3iKBr5c6/uTzaoB7r3CD/hJeO46xFqEqOc0Bod1oujs1WNrlErjCjuUla8Sff/3JC
nCdDaxb4a8HnBm1kp6QYeDAnwu+sFCeIIaYg/Wgkokvs2Y2957CcmCRNrM/lfjtXAyv6osNnyHio
mx64OQeED//is7irI9UiWjV6b4YEIQUULUlhLA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lKgpgIZ5oTQmuL8bPH/jhLd5oHLsU9ss3kSDYQ+xqDp9XqBitheXmzz0eFoo/aREO79ZE/VFAnN2
PKAMARxtXDW7jLWxbjCYS3EVIBefAaDkhmoyeBBFrJ1gmW3DiU7n0987Mv3D6+aKPK14C1h828BL
/oVWfXzXN95T+9+3RiR8ff+gbV7FSro5Hqo/lpL+s+shRTfHFV/jtREf1/Tq0qHfbWF7AH0ZiGUN
phFRWWGKwUXn6vLrlQ5k0n62UfJdZsVzoCQ9VEbHMPnvELmYMwTxSz1eHmPnJ1E/ToRpwh5RWLTC
2p7UpqqMhFoLMRj5C+C0Kue5Hf8Klm10mB0GrQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E0LkMsjK6RVWDWIVIrKmKKV0BY2wXrR+7EtRiSoP5cSUTaqGu2y1HMRimGo+hjGCNvkhjomq4fLP
OdpP2b/y1K4seWcpHMSKa10hDeHvBMj47mBVVnXYb00oMn87BNns0thdur80/NBf9qqnqMhkLRhl
f5ic0d1VvpItmnFrkh4=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yu/tBHCtu80T5YLEQcJFvzsX3arBNQeFBvz88K4l65OwTBApgKH2Ev4Pv0LYl9O7DQuDmOThg4qS
rIpvWUap8LN7GFKuP08BSJ7UOsOG1m6LhVxD7RF2j9abk4BDY3k1g0B3HsOSkWfQl4n3VMDLuwX+
VenWO88taiv945piuB1zpkoIUpxsO+b1DAnD99v+th/3vYRVFDq2teg2AaWOPKFr5BumM2qbRYW4
up/LDXhKEvMTVuMzphB2XUlYlpnJVqRuLZ1IR35y3EIUsUZXDVegx8BJswULNwG80NQc9/SwYBW3
xkpojnGTiUg1/oI4dQThQtYBq3v7ydVRShNPvg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aB5k9hasUxG7+3MbK32nkz2MSepsfrA9iboqLGwjdjKydXBqii5fghuf6OmcdDZrEViDmuwYQuUo
SFcRgxE6P7u/Ro/dAFIdhbbMIoOJT/NeVEXFygnk9W6plxvWNHljTJm96O7E+mx/JZLgv122/SWL
WL9fj5Lxhv7EiCa8hcAcdx9g1uNs2s1Au1YwA+0lrFMNVM5iZjQP3MQ9ARIlhSNIXZKZvKt6EwgW
yfF6awZwXOACiswawlZwt4WV59xPER3rCd2bNXcJPbhtt5G80BqGoM+qKYGHIOVRBqG0FJMpZLzm
Bb8JjjRXhceayoedM5HHBv/1yeXmwgzMyiJudQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oiRGHczAYhqnNufV35zDUrAyPWVNbE2CIqYIqdc2+7H2h5ozVAdGscwi01Cp+c20lPyMqwTWeMOS
OZFOjFccGif/1ehPJ/vB0Lo/Nrlgg/myIUfj3Nz4yGBVT9nWQXNkB+/U+zPpU9NsuwDgR327PE5J
o5npwb7RSCM0x8q8l70tvI4IZUSqx07ZmoGHMe3WT5gtMzlA+VUJ99g7M3qsKOJKy72Sfh0zdlA1
knsHQbjzc+dyvsrke8z29T5j7IQ10ggKQAABHWpEJN+O/3AaGIvDq5RtSnCZinAgL18ytNbQSyNV
TQzooPpiaueFQmNCkNGFTUMHShlcHTWnO5ShbQ==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k7jaAISLIucrHreMNA9bS5vDAKDLNSlmct8VQCwCtFl6abVDVMYbA1AEbizZSaC7VYKm6B1IHw3q
09XI0h4FHW2MCJEN8bYWIIjZ4sMM3I8dNqqu1PlaJaFSl5ewClyElA9KaR4+uNueKVFHnzSH58bB
GOShKiHP/9T+5+kvKbDY0PzyrR1yQcAeoksd6q7kdXV600w5XfiqbyDB1oG5xgzR/8kEdM0NEdf6
0J6LCvTHja0Cdoksf+7nJaQH7zrFM9ZbgetMzTRW6oFs9qWy7xeQJoBKQNiczkUcIYYGTycMXY0e
P41RIgR9TxM5LBjWbH0kSsBTWCblw8vUl4hPNw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55776)
`protect data_block
XKgqbB9kRcTqmwMUU7CFy+vUeJ2uSR0l9+kIhKRc3EiU927JfrErmWLF+0ez3kmlkY5nRWlaJC+l
Ou6Plus54iqHgCHjZhSqOLcdBoM5GVr12pteGHT0hOV05CdFiJkG5fzdKbIOv3ZjBlEUILKm8Jjd
zZ0KTyRHMQsfps3UPU+9anEucB4rHD5b9uJ8E8h8+oJvbNhs1pZ9tYR7wdlZJkt6oc0d05R8kas3
DA/gQmOgHNgyumBHu7/jgXG7GcYfMifAMV/XaLODa1elmeTZ4/Y1HOvGF7PRL0/PPqGoziTBrd9o
BGO3zIn/k5hyKjqvdusk0Qrqi4QKQCwQ5hClzmcvpHQGgfSARQ3AGm8310S3eKOK1fatVwkjbocr
dk9GeUDCSllLeBVDEh5XRhMh5KJv2H5wmPeiG3JS1QOBw19mzn3iyQlsll7ETPGJ552/h4vYIlZu
usn9nLhPCcUflDFDO/TwFsHfoewu/6K5nFIsX2JE+DhZfGUzS0H4YMtoaTTryMZqn6DPXIWEnI3z
HEIV71vIpvCjYCTYGA+XsltXA4vVVykbJSJBObB+Q3kjg2Dukqq73c6B0W5zFW4qet96CPHE2q4R
IgkPlHWEiBwHOHVmrRRBhzfPMGft+O9lNPTXp6oGjD2GMKuurP3Rvf/fH9PrcSn1PxAqI2AydQC4
0xv9R/JwZo5LApdj2vqKlS2B/dLZdRA5EcabREsTX3EkGP/RayftMZWhT83r3JGKctD66NiXW+Ei
V6sYUG1NgW0M5koepczHfj0Yv01MzBr63rHgaud3peYrZtNHeZnLoDgPXSyxo6IljhoVGj7hmsyu
31zOIfkxey/Pnx2+R0c2jibuYtAWs9Q6MPRGwN+xft3XMNHWuyGbyMQxQlP35TuyU1lumVvbXuAY
E0hzRg7CISPa14iuyJbUZOWQS/PRvXq6uBCjnDijjZxjKTW3LC083Z5ru1rSUSz0mmS0pcBIgi2W
hkPyxF8swJINzDQU10/0uTY2BYfJ+CgwsIoei2WEhJEIVbuG509zJ0hrZFFYM2f3Z0hSpJtt6A7O
pio/rW1ESsjm44d+spz7wx+ORXSdIn/zRYUKYTmoJlmWJzEAEY3yU9fTuE5v9mi6WEZ5dBHaXheU
RnEcfCIHWzVyNOKcqqRlRG5Mzc4L4bcDvurPEAg3B0X9hOfa4EjAU031VJttQyhBhBgRIJeer2uL
g7acoqz3rYJ5rprnKCZE8x8itJpK7tILkIo631gZ458Iw/BRTcHdiqel+I6cDoEKJYKVfxO2rStu
WA0npYFjYpqrcyqUDTDqRGLj8qNWc5uzat1S8PevCzaP++Rm5cqgFTTjODorzl2IpbgosuokLPGG
DI1N2kfxs213Ci9JPBxPnNXnyJVSc0dvcH3GsbI7xVe2EbrpxaJtenk26Z2+GSngSArmTFTakuUC
4Sw90VqcOkL71If94wtPu+VVB2B7MCJospXknMVoqFRIMyYzLRiO2u4Y/Rc5Nxf4QHyWNEkpdElh
WJp6BGWTLiNhjRE4h2N2EbHO2IOeXU/q/rR6LQpfxvCE4MHI6bRg/cevpWNrBZCxKIcGTSJGd6Y9
HwAvJKIxETHG0ilLsofIBFDhoSwnd+d+9XdqPiWydXfw16ajytVAWPuYlURcq+ducI6MDewXAA1F
XWrKG6eQcm7V5WDGVyPUl4U9IOyZ6tlkO7KTNCb2a2la+zYiHs/Uq0d+fTo+z0pVRVZFg0xozd4k
KXYeVaoZkPTe8X3quPNYVICkx9FYsRFPbGJh6462Hi6ZIqSmWZi3fkr5Z1QMO6GqYL9o82tlELtp
qW5av1x/gv9i5En1SFOY/XTxqCYnPRVXLRrP4MS7WrRVt7OXOriNu8OR5xCvj7JVoW3h/73lCHIn
KTAJzW5iu478kYucV7PUHI63FipgFza1C3hqEL3JZD/KGyyi9oQsH0YPXPF8Sg1BKmIDqN2lO6st
bD/r97fsh/u9xtOtOCAbpHpr/hpcDDjpmI1hexgX1xwUaoZg8ayN+7zztHudSPXolecd6yWBu7bk
VBh7iLb3c+ehi9OrIY79F7j2sNounWoweYON+nUboju5Ke98F6FSK1nQHm4M9n/eyftVv+2XU0R/
2csNeBhzbheUUiP+FJp4JtptgPGQEVORS5QFq2RtJdTalqpTjV8kTfhwJJ2q9W/ve3CjWZCdblYa
Of1r6851maNmU7ms9ydX5RnPkwpmZmzirCdpQn57zlmRDH3IdeVI97miI4/c9Dxxn+Cc8MTjMnd5
JuLsDT/lTKAupcAAD4Dj5T3ptzR5jdBDyaP4kFbGKJxaAkTxQPV2OxVt1LOj2LnhFTgbgvfWX0q1
8j0VlqDppY27ujaeTBYeh0s8gRcqzzMP+eIQ5pcKy4PSEdWa8BBqTcUNvwZGfPrre3e9VulgGzFb
wZatbzjk7xVfiIZKK28RldeE2KwBzfkFnfvA7sj7/0qMEuT29hGevt8D85J1xs6LkCN8fWxRRgGl
zQ8j5aGjLweIMfgLMtXXksankKZG425fKpfNwn+f9falnRBCPSoU8PH8zWjVHQu3fBzYW468o4TL
zuT8Kg10Jl5Z+XJy0eXkHU/eCaJob4ugw/QizMExXkYWTd5ksQmbf42CmgXym4ZLuqMyq4G4KZIR
ri8vrxua1Xo5HAA2GCnx8BTfuCU9pDIaGJW0ttV3Gm9/za7B+6qUwknsbPuas/9yRdDvrBlyPxxp
AzU9SL1PZxQr/DBerVPS83bAItpmq/NpqC4dopJuYeYXnPlv4UeYDFcsVzTU9wfJetLBkrtelU+6
dCw/JvPG4Fo6wcVP0lZA2abYWOSlLwLNIheVt6ZuGuo0BQql3SuuOYyHlBP+5vM/6fxVr54huT4m
DwSpuof733avawdsTaxdCDX5qTxTxgoh1bTRCemn8jaIe1TlSr91cWErbbz6ZJzJAhk/PBllWb8+
R2/1vZHHN/7VYntWB+Cno/N40RbFffQEeWWY3ZwjMt9Tgvejox4iE9iLi2uSg8KTs94EogL/IUec
lYo7lBNQpuPXv8YtLTnWblpp8VCOgPrs3F5EzgRhNH1qfzsrDi6ltklHFVKo6yOw5Nb77oN5acFL
gR+8eg0IYFqcSsRljdyHWPlX3Ljcbwziso3E+Dc9EUSgtYhP2X04FGbo7CNFzbld5DVEFX+r/zIB
nMk2RCmx3JfYg7uch/hO63Dc/aOEAME4bzjbQ/fvlkq4FkP/9VVnPsaguuKKQPt5DM5mvXnwgGEm
w25CztSc5BRX9NFfecoFKXKYuJ61oLSxCX1c/Ury2Y0sziEnTcxOL2tquafeUaVALj4lVaLZHB7J
q30qyvmqJI9c+qFDiR+lyjsRO9F+xIa+y2oxjvZn1VNwcGIUHkqOtbopi/xTDsbyyBl5wh3jYKT1
vGKX/5IZ48hrWne7rnhHTr7wS7b370IYLtBdSOgf58H7/dFWMqMwD5MCI7vcNX4x+M3r/rnz8L3h
dBPDVJ6xbKRm6/pVCTLYwCAH9ecCJlTNL7Kj74uky8U0J7lUZG2UaGdEVachmzgGwXUJ51PEC74O
E6AGDihH/Wu5l2slSwrSYtPdvNGldMocAYG0CZwCn4SjVslHzlVgnx33hEUcQLN1FgKgwZ9KqOl0
Rsou1KrOCKk61w/rFEsJg9II2u+EI2nyNYicmhIrULr//gT1ohbaEnVi9sQApBPDfAr2ly2lDGvf
XJT9xxzwR78c46dUYbS7pKfKViFREQ0An6HDDCHg5gRWsJyFHmor0VaQ9qGr+X43UnRrIoQs/c/8
I6DiQ+6vNlx4YxeX7viYG72Hth0yjxl93drodLlbCB9WWL1PwM6giIM52ygTA+j3wRYTgDas0Dim
dCA6Vpo85ubzLS0gIhvFGIdcty49tUx44+6jk784Yemkdn8dQ+1jhZdYelbDxJ47G3eLaDN5yMB0
0jI0lW/FC5Cb5PY8W2KcJTU5iVJa1FtB6FDh5fKU/mZuuqm/HtPi7d+TVJf6XBB1gRiiNwytFRAB
2nkvt6D/i8JNXFKkMwn28kyvNVF8ZZzOe+BSM3iq0x/jzKiaEBpUOrZnwA7fcYRD5icDWXli6YxZ
e95dy7xap8dPDLKvm4iY2qCEEPGG/wmmHFFUeSjQvQKaJSr8JAaJAQrcjLArDS3WLdHXhbsecLzN
X62eGjuN30jyPy50tVVBsLeXGb1CdNPCfyxqFk0AAgBrixJlv6v5agH0n4B4EmQegWkaOS9doU4d
pMdMTKmlypBdeL7QXkZA9zpMJp3UoeCAj9xrTD8MIG+fqeCNMJQlYM30DGcBQqfPgnyZiBVMZXGm
u47SCk4YKgwWddwSnZ3zLaXKe1VwjD8M02p9I6R9+qhUrCaRxxis6hw/wuP+HpMk8RMWDN/MW0cW
qtcj3dmnElNMg0d1sCRtfZdvWY2e3Bs/qE1Rw43c+3QXwo1ngMqu31khgDwhmUMrbh/8KuLAyqfq
ZGw68zD3rGjzAd8O1fWArdC+G1gm2kHYL4WoVlUVIM6Vy2JQdS6keozeQBsJx2rxXJvL1XGQhyaM
eZ/n+LlAmQ3ejCGpwBd94tDtGWZicfyhE9ZIxSrzP4+ED2wdLRaMckyHYCtgBxjpXCPkN3nQxAYq
GZTP8ECATYTPR6mHGZCaDtFGdZqIkRwheqvCBdpNZXtgCahLaq0yxBsskOqCqQRZaQX4B4L+2z/n
ZYivL9KM6nS+TcM7+ofGqUdpW3K3HZF9X1fgzGnC/qK5bCs++TjbGs4JuF4VmxL0Z5up0xFBnWHt
ozo3rRJFr+MXj2jb/IZzLxtFQWDDIIO9PNpTB4ULAQeBrmiAe0cgLEBIAFS22KOraqCI6wNUhANg
4SPhviigpWrP+rVr/9tIU2PE1DZZHa7+mJxoqv6NN7howLnDTtCfsyEpn2+8HuLq1VL/gRMwq7Yy
EgtfI3jz0pmlpYAPEMQs4bIpRI6C8Di/aHN91de/xQHfGTEtUKKZ335pZy3p2eZn/mXDTsS9d5DJ
xsPj09yKn/ed8+iP8DNFLmvGh0JEyF5XReXTFbkBcozybipJtmEsgKoZM0+HIDA/NMOFK9B0Gp/j
dSFZXGLqQBVt2J8p2ANSBwvqaxN6Rzq7gMn72JJl0j3PPcDtQdLQZyEul7S2Ge8AuwfRGlgj/66z
YFAiYVLnW52lBiKEVUpCBpU3yI6V1hBwO4gPppUQVh7y/B8Bz3l3oDJBPUbsE5d3UVR612NqQXkg
VA+XxW7Kbo+i5/8Ew1P6wdBzqZUSJptUJt3A57IttYUTLtd1bqQKaWh+IkLmrJsyIypK4oMTeZJq
75bhFf2QugIGY5FySbjPTB1DD7m8+AtnjQfcLCiAflDGrQ+w6zGPxwb/a5Cq6XXjuw/ffMb9u1u7
NLawJpVmFG77SXOkAWbnzgUgsYBHDOKn6971opnUBS9Y9XHTMDM9/LWEMtEcMDcZrtvXRWmI64Ll
cKF/vwbh2fkvdB3RyrfJTgKDlFnVUVCNPQHD7akDX6y1dyvb7Z7OhaFN8LvzjbFqrFuboSY9Ay8z
9YWbCesJVAU6AertBZ4srPFg/tPjVECQcFHN77FgBphmt6K6Bn7yfJ2amUoFrGD7ogzSd4OPw5zi
n2yiOqVIiWSwRyl7MOOPrSdvrx8cNub9Awj7yW+Hi2voluNl8KGzTEFftnmxJEpO1eqVAq7wGS7F
FPSTZAoIfhwKxiQTPSDKwekWSKp3oNFOz+ubu+R89Yb5tGKx2/pioAvnHVAqv8CtpGrqq1QvP1aY
goVzpqULZCn26gis3KDiMwGfId8h3mNFJkuh0i/0brpASrEleiBLPhajC3vFBXiJTy+DlbuzZw/9
nt6OENexy/8X54vb5lbyAgODDJAUcwl6QI44s2Virl700OmRx/c2gSyAJLGDQDWL56n8HfHgqNnn
EWEhqTWVkPxoIs/rPlKaJWN5G+k/9H+9VhmUvxuxjb2zvcPFm/m5TED4PRDjcddsJXy46GP222Dt
lUS9jeREVSK7SYjtsd5+AZJccsIIcl7Erkay5vGFQwpCjZ221fedmxKdqYb2kY75a+DLuR9SCoXu
fjNiLrHg/VhTYtOH9Xe+XsG4N9y/Ice9ZZPSCBl80GNuHSzZoi9plGpfEq4ocevZ5DkIyBRI0SfM
fX+dDeiny3C49tYqo1iJpiMYgkwrdzvhl/rIzeeE3ki3HAj0d5/Qq7ARmglNcm16IYflukY1wFlV
8j4mp8dvTiGOTuDvO86NsaEvJiP2WegK9757J7UbLGQpABvmXJn5FP7p87Wai6ps5mevAnGsBD7B
FALPR0lssTGFQ8F2EXsADRkFY3e4RAHx5fTkKx9+zisBE5dZDLNakOEHieTl4mMKgb5yQl8q99ob
DZuslNqtEksDr2MJ74YZLYsxOvxup0NTqcmccQE4BXaG1Yq6zu1aRzjwVCDBqML5oKah5CQh882x
4N+YQzdNmYtmYx6yWAB3uthW3u8inRuGBeev3oMqKznFj/UEWbVXe+bolHyz1OukUI/nIBTo+8hD
zl8+lpiUKcjEdLN5J/b/Z72ZBp6HAwhQ4ghG71CuW7HRMPq/2+j6bP+X+HsiQ7E7ZVmpv0YlN6ua
B9hsBOAJDmbCTQfU1hsJ9txSVeL9+ALcyinAE6UvU6jzMdSG8dRn9y6OhR5uB8/AT733rCBSxBg4
4WHe+siOa/B6Egc/OuPP6oJ0XTrUgGHhZ96mG4aizWBfors68tQuDE+pGXYcaNW/WU4QDAEXM7k9
riO000Y+di7A+5ftRPMLOX8/LUrRsurlKYa+yq3QP5WdnVLJdsRz3dqUmQPhbzxyiqxxdqaw/H3L
Y41vK9JII05y/iQY1qAlt4T18UC5GkcuEbED+uAhy5Q8b3gmDmdCgY7f+uq1QQSdn4DQ1gUFPK74
V5dZc5gRzNy1ZFWhoMFyUcnK24v//8EhejT3PlKLZc+ST0SC0Ls3CM2DeGaf1hK4wShaalCTUu+Z
EXxqiLzTu2TqRVllHy08h5tsRALp4nWMlHsvFotLWYwhjSZX36d9GaGX+Y0yoQKejEMsxMzSri1y
lfqTMiZNsKnt4tMlNS7tWvIPLQOtVdl/skCKUh7zNUgwoaRwLT4KkYaIdx6VeCAKDdNLuOk/M8sG
IiQsbuQIvkLkr9RchF26rDFN99Y/uyIh37pNOX+VPEqGf5hR0eL6mPNFiYVqAyy2whF44JfsZcDO
PqkQ1zjFpj5Pi23s+uAT+vwsgFsuV+e/eqgPBEVRUuWwnnhwu3a4apGbr2ef9EC/r4tC5T3M1pky
HRUXUfGCA53C6MZ3FhIFbC5QpDMH9BkXrVqjQGBdnTtoTZHYtRlwZnjdK+yAjw0HFubUAUTSio/x
A9lY4hgJ5NDIZ4OhrmN8+8I9R9DECN4EZClqgbpocXKQCo4TnjVPexW4GPjnk3wAo+0KHoDfIGmv
HSCpPmm+ECU6M+29l4oPGYoTncUxR0yZlYOtcUoKgitOrwQm2a9r4tUgFYEHZloYIB+JeN3wlzoz
jUcAcNkfX7z/v/DCpLdVIWlNbhP2P9eznVECmUa59xX8tL6vZ7KGk9rkZ+4TR9htgXe5/7jV6dMS
ZSi8AdZVDrqTGOp/RhXefclJOrMqEYsgoSPWdoLiNAWKdcEAbgJePV3QLZY+Ol6GOi6IyrS4SiRd
iPlONCcKAEsGgoLpYRovqu2uNSxbRwIirCgh4oDud4W7tF0EoC59wg85KnEImB/fRvhN56GuonLn
sOtcexbw5ebUWSUVL7O99bH/i0ie6ZUJR1QtmXmKRQmiEy5NTB3CTCjL/G96KEKmWvoURY6+0sgJ
yEBGDnvqf40yMveU1SR+/b/HBR77qec54GU1U8upVo+BMIQNz49Mxspe9/lro44HR0KzVzIy32By
4fI5y4j0X+7AXX/BsYSLRQBi5meLRJ+hENJi7YtiBcOo6Bck4Mjrz8y9woFuYG4c8hqRb+OzjE2y
yZQTaWkA/zyuVcZfUd7/pElva8tBnKcmZxZjgJWV7mQDGsugo8u65AwSw72MKjJzgp8VJnzR7/sy
iuiF5gvwa48eA4tOmiW5GMSghtlics5aMtsouZKusKVzBrODEAt6EyMAu6jQOvU9OnVHIPuB9d21
EydMue7aqrEcFJKXuk84q/yAnwY/C6bvnPLTARVzGbrR7QxU8VKjnav623fahAaRTf48Jb0QZAEW
eP+eNRB2IA5HP0ukF8uDqHWSeDT73jnfMWzAAkecrScuX7722zdQsbqKSldtZc7rQ0VR6smYJFfK
TIt/qOTLiIcskGk1H3BPKU+h8jGCuribeztn/9Q2D5oKdnyrKBSBhHLBkGZOcfbiVxj7wPJx4Hba
7tLIaVCQAmru6IgfkW6p7eq5D8M+gX3Phual6RwYwyE9E9vgxfFs98OrWyeW+vHjFQC0ib2aughQ
7JFRyobIwf8Gz30NVxYaBrPfSq1x3tGMVeK5ff0qIeVJJbkAbI1OrDOJDxSobimPKnNwlw6Omg48
HOILzfIK4shAzATTkbDuGZcGGY8JXFq/oQHfAGomgno6GBxBVTr9fwKc532zUPMH2X0yIUE2/t9d
x1iWU8IfzPjScV/Mh2V6VTN2a40tI9XREGMl+ZRHzqMvJdSFSXRIrUV7W28Fmu6A3pXmlmLiAmd4
qon9CztjBqgWMI9PAaApN+C5+rcjebkrlbHdpCPjsQYEg08mwFx67BL8jKSAjeAPcdLpZidWDVpS
hQUXKEomqOXYnOB7w+eCdpl86Dd0LONhNotbEym7RqXbmzCb0SGVwO3ltoIOah5KPMkMlb3cvS2E
OR8gGBpPk2HrzHRrCPZMAMqti+7YjWs6IRVL9m36fXN4NGO6RkpWBHLPWkky3p9brYzMKbUyn3D4
SmQ06JHWD2b5dh3N3Dqe+EU5rk7F/NdCO4DHd/6Pm+NoIKO+KL065Olaa7oHxFqYkFJiT0bKXKt7
7Xti6HxHCrI1NP8m2c9XzmbsTdnLmlD47etH3W6EUXQk2g605YJd1M3qApngYnZLVR0m/lBE2PbM
zdx4K1EXO+9BEJG8LGDx3BmV9NWArUXytPV2tWvALdFNmTjRd//IYvcovMKFsNsr9/o0xCOScPsb
/JbqtdpPYKLI9QVVCvXkRBJjFpkX91Za3XWLlLb9gIxMn5G49Y6WxEGZoCmDbOyreUm0K4B1JVhQ
0XVs3CqkRAHOQRMRZrhyNhFV1XUzQyz8LNK6LeRmfq5rSUGuzcGGYQRCHxlHmjRUOpfdSRH+1PC1
MRHGpWp+Qq8Lj6uLdwCXavHChbLox9DYHlXS7h4nSQ7gvpMtNsPaCPqtD9o3TesraUDfzMpHLCPR
r/yW5EhnlKGUkpdRYmycJHm1LEvI8n+6tE8igPP0AQeRk+Ospt+rQOTRs6mDPiZn17OL/XPcKKQi
AiKJeKEI/wjfFpxFX1Pj2/jBKYVHjKFynSb7VRAdPHhEfTGu7+2iM5OTlBy1E9+rf7YX5ZeOPoLo
tHk6Ggsl0DsrvqcQ+OFIJzv/Ls8RyVJ/Q+SYVJdb9w0E4Ce2JqRQacaPhaKu7E5V+rdEG2+l5pQl
FYQ+VbpVHT+WJYyHMrOBLziAr85ADFvsFZg86kz5EwWJIjL4kU7/vPY34H5837oONbMZK5zeHD0m
vlT1/r4pGaKBii2lADbYwsk4GH+AIggiT3uNL27tD0WiM3wckQROXRfxBjlyg2ZGHQw+ZYnS3+TG
C9oX3SPQG5t4xn++vsr34tfUyAEHKBsfpP+N7JT6h3fNoep59d9djt19Uw6y2E9JHPvx0Y0PY56K
zNJvb7R8NUNJFib1VuF8C2UOBUiQSaBZQcpfigzdLnV5N7K9saTLMknC7elSTtFqdlpHMyr/3K0n
NHcjMyIpWHwHS2sXoydUxsI1ksnkPK7zPXK1h7GxWVxLC03ctkN2zxyBgPty6epCgSLYIJyO2wKP
k4CvR0rzkNbivz4Ek/C8iydNBiMgoFm7zSEoybJ9kNviaUi5k/y82rG4PqMADoVEhJmEFS1H9AzZ
p30kPBLGqszD4JaBXT9MGRBFKqkdvawKHJs706HrBQzE2oWbWImskolsUB1fmsKknEjQ/aVdg717
uuVUXNbP3MtsxifwApuKcG5LMWTIKuzQE7A1rlgolpv+Qhlt7eoNChr+yWxdebD0BRKqPNAl1Kxn
m+Q+Of26hBEHd4Y2wWEamMdVirMql6fW6Ci/N1bMHHG48szwVMqttH/9e87RjpKHe59B6D3UdBbT
H+OetewyGJkorgP61M4tHyLHRT8fKtf7eBkgpOVSF1we51ntUA7csNdXjRZ/hRfBYNfuyXT5S+x2
dWCFPQciGSR/CYo/TtACUtRsdYvjcFOXGUpK57yWJFwcUF7L+yiHWN7JrbxTGAcQGrLPsRmr5V/A
bU7gwD4yoBRSJVfDwBW0yMF76ptimjKYJG0N6We1ZXZoBD6Po1xD/DnuiZJKMURuZq3UwbeXEAhv
yovBQWL5Oqf9YqecfhhtPdcIxVIbfZ84xBq2IIbtgv7Go2b9L18AjfUwGZ6tX3xSY2LLINUB5Pi9
PAHWDSEQbyktml4f4UX8r/ozWZd5fUVfYqgWUnXND/OsEU3woG9O3i9F+CMoJfVUVrsmNxgYW6yg
XixvZRs7GdnYJ7FwuWEFxdjgTNEGtOsvugEYemH3iT76GqFMKGxr0kbW5xGfFP3kNKDGGn9XV1NK
lD2TsqooKGrEVLPg3Fqq5521jMqZwYNzA6PLp/hkTWBeqeTfrJs3w7ASYBDRpGWaMJJgo4yvlRa8
oeo3Czk4W8UwxAzJH42PgK4nGS+BOtpu7el/AHWwSJxq7zVP6xuB5MwRnTC71WNn0y+gsiCdB5KA
r6k78vBO8mBtEn40qFFPVfz3I3j9T0mkFLlb2ER+l0i7AsPpUkdP8pQKZUs5fWwsAmkBpMOdNI+O
KXqjkFKq2gYCm7ZvSwyhjTv42cMrKPTKnGAEeJiEoO72RtEzFiQJ/BzTIPXN9Iakmp7muOqlTUgo
Z3zm0hZQv09lBnrrpWQheosrUkGR5/6CTLaDoAOboVZEdk2694BjALdbkhXYLx3eFR/kYvOATiND
0rRn6u2tW/N2Z+pa15oheVUA6562/K1ABoWQdw9XWdos9SFmQidgZlRZJEYsvMEufMlMauU2Ipbl
yUn15DY/829cEMJx5epTL2HaDK5tgf9uTph34jDh7406V78c8d4b0DMZHkSRtBMSeJQtb90797bB
O3ePTqI9uFmKKhm8byQwoCKRAQQaWhcshxrJeGRN75S3LhoDk4rxj7d/LySIeym/sVOWZ9Q/x3xe
w4Z/Lm67CEKvpa68KENouA+gEbgDAvfKIsMUkTNRpwTs1W4KMoobV5wiYEXD/GoTTSxpqNQEU9VV
6E1XMEa8heYLxGUngjtqU0wiUscRtaG+aXTD6nRJXMyuWH9hkIlz1txfyPdfj5YV7nx30nvo3d5B
O0kfVsc5paApUvOQ+scpFW1VFy/jMMZBqF1OTrjJA6gEw9dAM5C3NUT8rYPRz2fi1M7hsjQMAeMW
vIh2kW2mRaXyupnNwwN2Cm9U10Z6rIkQ9VBylwZQ0BvYBhVlJlmszVFGi7jFOKj8jWhPFeD9NL0o
2SNxJ+PV8bj7FLqQx0axQ5yvlBMCy6677V5Ya5SpkdSns6zyvpBOxIDxOUhzfrkK9BSpE9xZDo1D
bUl6aK3/iP9ndUn9WHs1ovxigoK8EJnqnQGidSnPHds5IA4EwkIWPGS3WVsXYZfYWS/V4itsgHN2
1p3YfAmMfKpe5/uOaANezURHjZMU7v+fmdH69KzS6RBNExvRwOoTfjwL4WVYadn3QueoBUHIBOmr
YyGHdJhPcvGp46yAoCM0GNfyEO2N2L0VZOVru1Xy/hRHEbv2GT9uwMgX8v7M+DzQ+qVXMwrDwOmg
qqbnJYt5dI5a13foT3hb0o4iuTGzKTv+W92ECFrJrGR7WOWg/I0ofYpxAQRm3SCcxsdRzc6gyKOg
uaHmRM+KdYUJMtDIoq5cRG14da66eutAXRQV9/uSvmUOShnORopk3TlSmYYgtaZMOciAx2HxOkp3
zv8oWGFsqKLVRXkRlWbqaaPiz7wiO/QTDWRuA5tYdmrNY5p9vO7vWfG4b79B5cJRZ/aTqTyLBbPF
QG7UAOj5P1IS9VPsIq1ky7AqqqeqGDAELA9oGzBtaKMP17XAlDa+vmm8MMuGSnnR/TYr3EymOlMr
0L4yatK9fHkQyVqi86khLhUfHFvLiDEp4HekGewdq8G1ZCGZeCWFlHP3rOv/KlcZcf2gCVRTtHlG
7VjJFZu70PogeHaGSUvZFfkRdweDsaCiZWbj9sRGIjP2w5h7iVLtdz5BqWs/6C6nNhnpsix6DLLM
ce107EW0pYAT7YfPQmKWHd3laCdMDi/bfB2/1XGU0IaxU786GDFBTuo7vRjWy7DZOXsPivDP8+lf
GK1fCZlNI709mml2Z0vk6V72PfAmVYpbE/ONZBSWtsEffUhvZwZtHXmfv5JGI9vCw75AAFc13eko
os6Xy8oDGf9B/B4zP8qEkjCO1gS4T7bO0FDhCncS0vhVTwKFWPCvpTNeVghsxcKxj1iviUA4EQvR
tjcuc05Ua8Nquw7lFBwVp/4IMo+ZN08cPli+YuO7KHTsLzlB7NiJeoeXeetLQwWHkiX3uLPhc5U0
nFebVSOt7nlkanFhRYg8ojXAqLHH2ZwAzPS2j2FtGnOOTyYPHbgJ+g2WEzrKtUSSleqzc2zR2YkT
dPQtV/P21ECZSEWv5oBuT5c6rUL3ZOQ+7ljxhI1pB4vftGQjLMNwRKnKT80ZRE7p2U61bUoAD498
clJCVHPsdNkTSJJmdHff0AooKu9/hp8NxKePlE8EiUgyEelKZzoQXbHzrpCvEJRmi5kEWk9mjMWc
cVjq/79lUKrdxf2xrO2PgBOmy8KT8zgBxDxGKutq5vMJZaiUWXI74pDCgkisvIHMiLarhIn2zwsJ
n7zG/5V3kip3FREu9hY+zAYVE9iSUo7hIAzBoYgRMNoUmUuAfgqz+23GV6tQopcluR26ZOlDN8n7
ZVrimYz6do3NgSTf+maBJcZOhROzK3SLF8WQF7VBlqC0Pv2X99cMNL7vOlCbn6yDUIBv11H2D+I3
bnpeJgxtq20Mvmg2YpmEgUwnkvx8W5LBd/9ldpuSP1iEvUHKMLTBq7HNzhvGrAVZoBjEM0Etsw3l
YX+bAXcaseh54Uz0BtGSS8TcWKks0LMj4DpPqD8KfNVMDceTf2EzmAC/9tp5berl4F4UnHkIrqSQ
z+o5mXm2/JBZ6FOpKN10cFOYBPQW/rzM+xyHEK2soB6DaetBpsSltEHHs7tHpkaMyKEoY4ufHAcX
mC2NoQOAusOxk3j0OHO8Dl9vuVpnJZ0G+SMPh1w3pj//vxwfN8MnjOWdr6+FLvWhIbeeAntoU4Xm
iKOqC6ZrZDDWWgXN9KrLwFycC2Cu1S8rws67pKNX/xW4G4mKkfX3ctLT/iJerUlpeJaGVI69hZMW
281scVq3AXbN+AMHoz66P/CAZyaNMRnMHlS4ZbTEATOn1QEqUxeb6yqRkLm9ZcMfp5l12EUXuP71
rhUeEKkWFdMjULIIOXKelJiYA9KO3dMDtMAb+B6agf9+4BoOadW46erUxP3adEH5PqiDquhxArZO
Ov7juZxanjEeEGNjP5f9JkjyMxbUYSYqIbk6+YLxJh/u8vLYXlh0toEYiWd1cT02l1zu9jmuh0ko
Bhq/GTJ7LNeuvL+mRdVmeZUHmUcLyeSuntvY8UY+iTTdp6c4BcuaghxrE1Z4oyJhTzmN9GWAIUsZ
E/fOXs/E7lfSmRWK/f/+yussrt8J+mFqRH91OYq8ocOXaNmpTd1Wuk/QSTgrAdP3P79bqIrQ0IlB
XMA+DJF4vR4Sc+SayDIQLVm1QZ9KlnAQmPV+/PzMdDLehKhhwVmnbAbUM01DgjEYAlPUQFEY7vyX
JCDNj33UF7g/pixny3rKytvxI6xyn0ukiziMzXfnRnTTyXjudi/+Vjfnoe4zpPXxW7uhG2qvbSsu
cAOj3g13BTZyy1aFr1ov1Um0wxrAT56uQMdGEkOZgivGpdZH5dZhJmxoHFe91Afg3ywZG5ufhdnd
NAz5RBBpZJzvTs9iOdWUpvEW0gaiXnqW7Y1rcGES4MyMYDyfQq4JDVVtP1eCaDxcLkCQFHXrX4Hl
4ILjBnQXQi79IxBi75gp9A/0fanB/Kmc61xb909hd8WS7JTuZwwdyebj2uibUOJ8eJ2z+0zg+o04
/GQtpoOBd2o5lAxGlh1V/+5VqFZ3Wv7XSKqMyApI5NeEVNmpD2DDc7MBs6AfUYbB/eSV2sOFjpvo
qCnEfB0ZhBcWw9P02AbMtwV1RFsU8y8awfrW+ZtiUHwakqNUNRpUiUxew4UzS3YNfkIRnnyEOxOA
Xo/umOrNvehMS7AADU9Fs7nhxSrn8TkxqBIGVHIwURDyDfirTsWbcR+aNt1P334HBWyrOJdIoAwx
zPjSsBqEWlhHESs9FLK/tzAU2iGb0IH2F7ZUiGspzA7SEijRWrqqHhFC8ub5sNC3dGAn+yVfFr/O
xCc5h7+sGdYXdtfxtxTQoLWESMuG7u16hiRwYwPuWSn8Sit7bKLLPVdMAftqHJfwf4C5+IZSuuzC
mPvCrsZmvYSvZCQ3YeN+EcqXX3tDc9tuRaEKDLswjSGoC0E+raTl8dasdWrLFMCASFxH6sdg4KM8
8wMuRJyzkEJPr6Bc7RsIJIb3ggEiFQVQ9pIz6zK9yusJYiCyP9CJ5n5u1JC2M61wwYlCeF5fSF8A
3WvivRkkaX3EwF5Uragi2P4TAeNvKJ+mQ1MPDyFHj0+x4Ru06OP0hPYBPKPCGFYAi4aurCKEcI9N
mXxQgjFks62mUYnshSsvKyniUh5HOxBufQ+VOjth7jrO74+SQDmrpCnomGgIYlHEMFR+AkQEc/Rv
Ha3RJe7zvdEE/8sGWvteic5zanQhAae62UgHRRMoKiSSiRTQqMaAWozzLXTLRwb5/NcOrNvNHqxy
0Fzg1qsm3y0uQ6BP5C9+M6IO3EHaPcfJnz67Fet6Bj8US9P1c8F1pOvsVBBHkgn8FzmXgp+OxzCY
/DE8+X2Qthbia47vkTt7WBauVXmMPdVFO5qGR2ZdCzirQd3rIqQvdmVwmnO3WANNrQS+7kPnGkaQ
Z7amQSgu0QltP+Xj84rzsMCHWDCyqmZS8XUJTBA1b3+TxQa2+17VpTz7LQ6MtAYOKmtRQ+tgkj8x
dQCnUGGxwKRze40PI0GGoftkpd6BHXDYY5VhJNzEG6NzgK2Zz437vrPkh7sVA470SnOb8CVg8hmN
z7wxMF8Q2bcLnh00R9hBeuBYiA6jug5GkkcD4fut4UPeID2c73IlYrC4+GZRBDgU8wW4CQN6HWdc
qeN8XjHjPQocSBYZablpddW9auFy4g1zl3mEQU0r6A8f9ZQ9doFVCcTVOQ0ZFoea30vK5LMZ7mOH
eJ8KnsYIV8oTRLl3f8RHx+q5/IENd8ivjs6haGCMvWKAXSTP3tt8pjF2/CiRQABnlDBpEK+VsnJj
vOpf0r3BoSjjO/r4i6EY3atvsQcG+rxxIyFVHMeilm7380Om2I5SrjYcVTyXdDPGrduGRjEdun/i
itSr0Gc2LHQhxPs0IE/AwmMJwPKmCZCBQGdFgRMNnxjTsjPYjoQFmWe1v34a29GGyUFGXnWE4wy9
nMdGz03vjzqr5oWcjzLw34eewLZLMgzdbM6N1cW/yLncQPv5/rU1qWdjxf75w++MOP1sWIE/kVhf
EpQhDa3xAunLDlUd0jasN2kJ2OqFlfzaV6xuq/HZzs/kIV0fQxX3tre2Ng89VPRGTcPYxQFsqqmp
laDLpWx8c8izxAlRLltSNKhTaQdSbSmTxlkfpQYvCRQxZ5Cun3FWqpdxgJjNNuyzseM7Z20POiqb
8RqCDOEk8rw5piKBhfXuZx2Zh4Lu1BGylILyBd1XhGViDoA4oCJpKlyLtxDpHKfsFKZP0WD9V3Hy
9Idm+bJxRyHjwbfjbDAVV4pueQ5Hho0kTDij2UQOVYST5ciyIU4631tMbwrtASQNNhO9O5MPJxwv
YvkkjV7FeI0AogWojxcvVKpVtYArMP2ZIUZBRBZfBdTgZRkWzMHMg6CNOUuCeRxLFsVrzYhjkQbs
bOTO/KeZMQZRhjNSQPCSCEu3zT7+EW1+jnIxsv22zZk5eMCHw0sDE/m4uu1SXU8pTNpulvr0/ORv
X/J5DRi1ZtlUAbe9dqh8l9b35YwXRFWMmq9+9dcr7xc50uBp4gF879yWcK+azxBOMvO4mphSeIHL
sb7VZ31CTN4WUnMwnUtMqlQCdZ+Mpvp5bGaUSqwyBvkqSj7ctlHmDiHX/8DKuxTuALD4UKa3Hhnl
3tqHKTqwWFCWzpZLAZBifJ1T3HF+B3s7s1Cg/x0G5TDnhO21GA+W+6TE32HwKfS8DA2FmPhy6P7U
nQTUvlffYirxZ0JqmWug3K4DNSRjt9O3+3c5ccQ+W/Jq5za1XaKGJuT1cqL5ngBPkvxdSg4qHd6s
VSVv7hiog8Cvz6IAjJfdoBpcoIICfrq5xBWru0Oh9ZgF19gDUHg6Pj70ktwO6E1fPR0PLcUhFDFv
8GLTh2ZgeZUfhYDOqPhn5RWgR4Q+2e5ZfuXslmDOOhYRUVVZfWrO/q7n4f34Zhh9BAhuaDzbuVRS
IEVKEGPh1zpdLrYwfy4GKgC2TI5jKWhCflIuYOSgJlEhL0UjhXn2DWv94T/kv3foIseTS0HX6teE
meeXx1nNqYNCyBuEDiGLHiPY9VH23b2O8khgUyhb4Yzn9dVke93oeFwTM6u62KtTEaP/3tl0XNZk
/0HQdb93TUsTYsWXjcZCDdwAHVJbcYPl7O1tmq8U+8OEycYOca3fsmJayqZrcF3zBl7HDw75gWQI
znvJ4KBXZRHkMQxq9yXiWKDXc97TNVXH9M13ha0uXgW8FnLkgpgcfZBFF87x2U0hpe4kjorXBYy+
AkalvBx0w9UtOkaXbOsTtjvjc+7ZgTMkuWOGOkcUnI0C5HllUiMxiIAx99diEt2cRhubKpqL+EVS
7JlAJRTnBuVyOWl3Ns40SR0ROyqYB5YTYXNryi6xlurvznYdg1ihuSATzxSSfuTTaQ4/rvD5xw1C
KsS/jBLD0zj2Mr3tSBbt2Vh830d1SEF7fGcUfwO+dpgRgALrYheudIrEc80heSyJe+UAuDOPktYl
enmizy/Y8MYEfIPFWysicXiIcVvsyoV8a+0KhJivEMfMqVZ0aC1hjPhVXgaC6ykXCg9+XUrEmKI3
5GOnsU8n/JB91jsXxzqbNSUC+XKHq1B4jFIG4UBiP+isMIFOIFOvgx3GuvxSfxmV4wnA7vs8ob83
8jHFlotLVzGC2uWDEeJGy7Gn0h7b9LRhcqClFlRnJmUGJdDAFzsHhGjMlV8tvpaUGHzRc/4t8kj/
mdU4t0hf2M5ifl1TOPr9n+8Wc351LGBliNzbq4XzgZqAIcPbJpU0mutnHqEFL0GuqvPtK6CMLK6N
1rWrtaNG+RvFQNxRkBMpxQz4uJIDj/ezlxvE/oRVYy65Kf3DBSZ4YHgx3f8+c7j0ES9lbxm5T28I
xkBGx32LR5L4ODg7Qh/XRzi7A9lmoC+U18EplBmx8TttDzWm7V2x/X8whBh3K72gI7mR2u83EF9x
OYK6me6lHwYk7iPRhW9kt5Q5bFANSPR8WUj6U7t7OpBixCLwLosUXe0SY5aBSjxklfCMeahSEPKl
tYGQWt+naQODD8ENvQlxSd8jkJ2F2iEOcFCRz1TV7uOWi4uCgNBDvil9OXgzaS41Mr2LortTHc9B
OVWjoOHQJ058bZW1D4+3E3Bx7BNbsh32LTfI9CKxegkTxujtNJoDf3yvJevZhrpXvLoUiUQD8uyK
liLWp/T/xFMk8J1s8cvb86mFr8l1SPoHmS0FEgngbYIGgVC7DTW77WrDQ9Zp+yq4XXxOoP9GnQFa
zZseQzpQF6KGTsSJn0cVVhKRh/aWSFmUWG3Kc6VhEGH+4BYfbfIdF7obPt34Vy2CRSgBHnllQWVQ
RdNu0JYRfuhToy6oe7qNIfQkA9iI0Uok1Rw/YyfzcbO0lYwOCJplRvCEuTrZDwbzSr/fxz5OVJWa
HXFPEgRhulZNN3w4RnjEQr+kbwaRQBuiUJHc97tMUojSxn+qXD0NDLtLAPtoBdkkvuoparJv4SXm
gFW8+JvKJ15uBTWJfT8he40hZtOr2vqzB+ggYUO+f9PIEAh8l4Yn/Og+ZZAiJkUAdfkb0QAi3pmW
/RCjDresfjYeBhv8NrRY16bG/S76MpfSAbHn/mPf2BNrs0voz3qv173ezvgVF/WkqKbH2HKAfRCD
2FF9meg80yJQJKuC63chLFMSrETL5TjYSAbcGZ/uKsuqJTLUAPwxhXJejfVnGA/481YiuAfrG9Ag
MTtTov8lW4Vl7zY9doAD0UcVj+kruIs3IQvwKsPhvWa/NZthfELiRxzUbzbX/STfz/RNEPdrRKN+
PJm2Gd9anOGXN5Ms0r/PdxOc3Up+6jvsvCxHS3+n6CC/LCqxtBDtsbhoZn8xbw688SGZvsAptA6L
ImPJvXhhtOvVq2+HfVhpkLtt4IxQzHhxBNuPLqEtcW8DmmC+IWkGL1P+k9YN9zo00t0+wzkI05ZC
cUIrRY0/CWYwbj2GeKsW3mWcOF09ABvqCusQFeOAGnCEcdYrjchucmTsNR+T62EnLfKdRIanxIgM
ZttmV3Eh6viAOdf6LuwydFlsCS/4mr+WAp9c5uM/1DPLSt1KftYjpjjJn8YCLHeV0Kgm0FePyyzT
iFIwIkkC2xJUcTJE11ezGQeM/z1pJF23Q7RloZSstX8oVXTZQZQ+DIZG8gYOw+rm6e3RnnmcUB0G
eEuZI5mTKk/daAs/O+G4uzH5rKaO1isR4g/Vqf1iH8GE+OSY06fzAW0wqD5CZBATXrVod1ALM9Kv
clL0T/pqnwFOxfb1A71eArgmzHWz5WkVN1ozgTYsdQ5epzgG+tZHQLFTo6b5BJupo0ZyQ/xMVueo
ovlwipQpPuW4uT2a6j/9nnZunsccx/VO6JfcnKYyahsSMy9mQmorS9+X4p0PShHIWGQHYbZJ5pxv
c6jnzG0S3VtaptF6BinFuStrTqByNL36FnqYU5EdN80ceguEszrWmaBbW3fTC3nXCtO5TP6saoyP
NtYS7i1NgwEkS1S9VTz/Sz2Ijs2EMznZiopUn5qurKbXArRJ7OTAf/Ttc8wDjOGt4Qna348lcN/U
yCvLO8OXwTgu4T+zoP3Qv05XERqeHbNL+B3PhKoaQNS0mhx1iEPk+riPrGwJXc4B+jt8FnoRp3nQ
nEOrKHiFvdsBFstLYEzhXqLSoCCAmyvtjVgjoCoJPUZMn5ra63EwpvPrLAP8z0BZ5pW/NzV9KReX
MKN5BIt/D4Ps6PhoHxpjVRRNIILeN1MdnHhSS2pWFgQ8nsNmtFxCLt8KuOdTiQc4Oo3wLDfzpifl
Enyu6ek+p46xK5mEkV2fwuSTucFkSW7it9bAHea85AH6WJw3wqGUj6ZWIqQ+2jMap2MfqrRPzYyy
jINgt0Ek9my0QuTbA6mpGty1Y2XiECRJSsI/kbS3UuaWklzvifTu1leLqQvot5aYVj6EW81CPXJH
nNbmU5szTRWli+Sa4FmslYdbZh02ST8S380PSVAHhu+wsTanIsQGRUOIQ1K4eEajws+b/uULVoG5
2uy6YtQnQ4kw2jpUJVAiNIEix0Tq5ULEgAMErfOpHxW6MrR6s/2/++27LB28aI5iceeH+4NfdPZ/
G6MDGHFIHVj+jQiCOoLzcemiTz6+n6uVxlP3+wUWaBAgEyrL7EduEmhcF3FvkQbdDtLzH8EOdIk2
96azfNC0sNHPdElmKez8Ir0UR374/rqTGgmbeEso/mLfp0v6Sp69txGCY/CPklMt1mXacJ234aps
7w3fUwUDhc76jqwYhuJnk5MJboJl4dhQJ6ndweQ3rrevVoIJlWQHFqDoUDCgldmDcqx/RvJ23l/c
MTEw4vl20XOxhzBLqzqRcXa8GhNI34Qpp5lzdgKJZWjszJXE71PYDtxa6otSL4TIzmLyxYs6D8GB
D3vAeNE1yY1g4GDr+bn3LV64axZu3677gB48PveC9AjWTJN2cvb7tdJKg4nmWvUPT5ZumwSnrE2M
FiLB7CVBjPLUZocqXGkdFtfezy9EXqQ0JIicwdtt4uVvyXiymlwHWnbGgzphGB6J2CNQOIQ6DFoY
X8Bina6pUMykP/ZHlHWeFm74rnpGBcBkVYJku06bUawRzTvZqCVXnLy3UkplCw9BwKYdx6zDuOM6
JpGgH9gLAMb7k0fHp+1U49HOthCEtW+un1ijFCdGWxgiHy++y9IbwcVEs/xDn8fRLlUeGaeZ1VBm
KkHxHzFPS1UBpigZFO+okeUuGBIbwOaVQyaL9X7sjB8MggQgcd5hQWw963lxuQ+z520lRkp9IEBB
DNkkWrSPXLFpKhESF5VT6cVbgT9STJiH6ktdtYjQ/ceMJWGpUCM2xDj0unza62MIkb1ligR7A/BR
wetdGSCNSk8u+en3hJURW1VPvj6Rn+jFnSmPjcThryzwhETFUTyHr9moPnTPoufSKXMjEzbQEHky
YzFHtwbayyyTregKGmkam2rxuZ39iRtO7brxH70y1MwCT+JJ9q8CNhMH0+P2KafZz/J3XY1Ct8Nz
01uC94202EPeFmChGQaXy+fVG3Dpk5d2UszgTmXgA98HeMKOIqsdixO/b5CUho78vpIEwSf1EANo
kp4DkQD63txsAlbXmkHjEpC1rV8WEORgkOTxJ8TPSyzwu2jH1Js70OrfzEELarnZL0RglY63tDTG
ll/Y69NhF+0mQxPzC0ANAiVSTyfccHteEEdH+OZbewcHtYGgTG+9lh8acXX/ulpo+HHb9Pt73N/+
SxBlKwTzvB9BoKHT4ihILExno8oVZLXI30DHeQIh0QPQEnzqfkq/7QWx0r/DJmzg0EPeTqu09QnX
mx1Pc47xqcLjCHvFJv9EixsEO8Mps6A59TAcfr4uY1g1THYE5RcXvk1zcXEb0ENKBD3e9O+8vjmS
VqWWKH1U21PUOV3RMrN8xlHItagts81MXbLL5BKEeW1D81XAtt/0hB8/4xoXBsHVEtLvGuqjT82p
Keu9sm13PwbMpal1CbEducKqO6vf7tLUoBN1msvqvlZxacexzzSGfpm9K8rNd8Zr9pS148tEoDsN
YWk+u+f2tBOZdOFWG4o3RboQ0skbSN+XhaqEcgW3RjBPe/mAIESUU7Lj8UzAja/t2VaLv/kJDzex
G8HxXjJkbwo38aEIDxLbM0ARd9bwYul/x+Fxtj4RQ4Re3U2L6Kh195v2MpPQEEUm1100GH496wPT
OfS6JPjDw+kGgfJT577fBI/H7Rj6G4gzmCknlwnhICuN+hVvFymnua/BUsboqhqaTvkBC+1eT5hv
RgCYXD5A1Vmz0XcywTIgrOGEQHzVOEKeo4IDH9i+IerWjL8EYIC0EzUDXDtIgKWSWIvHzW3xTwCN
OIRRvADNXsDKtArqbfVWijNQWVaRKs1veNi3VYJJHe9cAw/iq/eW9posIagxkfQwT7yx2JDAqXq+
ijCNXk19kf75bieHurktboT6DZyn5ZMMAj8ZbSjz0T7KsMchfjNBE6iF6S1u0ssw2XSAHlUjRvtZ
iUlyhML9EhREjcghdOB1BLdPNOuCvH4lDG48c+THikVQ18YB2mwTM/+VdLQbi/GZpxQ2TIz87liP
JABn30LubQz++ItxQ9ANDf/aTK95tphARvLzjdFzbgr0WRA4G+CKahpYm6bkWrpDEcGGsIPRZw7a
NcEmDPd3fSOmqmHIcsoS8h56x8Sj1hFYHpyR/3iuk7zyOYbD55n7/df8u8bukTXn6PHyo7wtRX+o
WZxHr/zt2WpH5iibmGywplXeVXxLJjCPvVIrWBY3x6rGOPLDeGZma3LBHn07gx3wDIdy6XwbyOXc
24TlnowV6CZBJIJsqALWYkdF2Dh/CNzQ/oDHnojN3d+Q6ZBzC4iOEmWJ2PFsIwTZaiZdK6moNSFG
tKoZOBadoesibfvRHSjul+ebSrasa6ZhTBcvySRhhF+OQRMk0vo42qUoBnhQqW4QlzJrhtMjPOU4
WQBJsOCRNGQ92/tfe6sW88CEP8ppXhOc8KGAtKQhTae6Cl2eJQyYXMjH+JZyr6CQUizxAj23KPMk
5Zpy/tQ93Wjh/kL2oWVL4W3a/lUxIX0L9l+RpzP6VnjvPYt1Ka3ruN/HRrEMupglTF4CSnprx6py
sF9Is2LyFqKeNEleepAHnSmyXOVboYwUzzVXml2XZUpl4tpGdO8Iy79hHa20mlB1/7n7LFkKLHP5
gopVBbCGt4VGoLjmpd2kA8+hZ1NFVlRkyQMWwglEKbdlT4ofWIkQ3N29rxEDfiNzlw/wiMPvAspi
V371CXzpyg0czM6ohrMHy8Jfi84SNOXyZ/Fm/+bOMmwKRIaRJ7cWobZKd3A4rAv5cO5XXHEAwzA9
1xEZ+CCU1y/rgfhQ7NY4xNqg9Zez6HqrCFvVUF8lX7MFpsq7/qXs0IxHUkFKNzH/sFSx8uM/Ud52
H2OLPEGxgZ/aZzLhiXTk/m0hG5PJZ8hwqLRRRxepMLpQONn8oPE6sk2rWltHPuwqUL3VX9qqQAzL
HijDTYVjjjPsGEPlbJIEQ6MKqgvnKNN3yvE/9Qlr4G5Bijr5XmvZfN28t+DDtFrSJvbb7A0no8oh
qrcQLe4JUtSRdul8krFMdapw0dbIDO3Js2vf1qV08lZcIx+9aHrdTjfzi9AYouEQbWToers2bSSP
QIy8sEJ5k7msEbcg6ZHSAMerdbQSz5fi5MZLAUf89vy/7VTsyJM8Hd+nQT52vbYenWbt8R9Q2CJM
Ze0syykOoqN3cBEB5WA+YsWNyHS+JxG3U12ufZtv9S8ObWg4aIOn6/gwo321pRDSNqA8jNRpidx8
N63kVRIlBbM86zJFGJQuPWtkXpRvzTJYnSoh7Q3k+3QlKTuImYTgPjdzJ328iHRHHK5DNOvd0Rq/
bXZ28eSLIXGTu7WyGnpkJ717KFcccUNVcB1noLLsQhG14mc+lKJreEzqK02zILYSlBJnCJAtCWsV
CX7NFz/q+uV5PYHmpVoORkEBKr2GLzOwpH9+16CfdLTMB9hRzhc6/P8hM8N6zs0WYoXV2p+ZPeWG
p/MkVI+iy2Pa5IGSRktt3Mx4U+JiKtij8qD48f85gzVByBjMBMji5YstKQbm7PmaHmGNHLYm6nmj
cT1qbATdFRCSU2y6K+9YfSATYbTKYirryTNd847Oi/4Uf4TI/tgg13rjJJXYMZsoN89j/eLzTcIT
eWkCO4M+43+ndE5KbCwbj2sU9ExQ3zM4Lkgnscth0xUP2lUSXPv504bks/jqfVrC0C07YMa84WbL
jpQgT8p1O1zSB9pr63h8RWCi1UMxGk5Wx3/cTpcDGvzdDTl7m82pCT90NqROOH0bqF/v58oEdQi+
qWTssskJAQicpJ1FFP0UAhyakUWxtDA8ksugL2dkrAlYGN+79C2MStZNZhI6BQ8mUpN+svhj4km1
f5wXaZF8Plg+tabcwuS0QWW2dvL0w8S/rY4CpgiCECJvQqlJxg7ku8YeQTQFShCQEPEWgvF4e5Te
kb16ESeFewCetpD848GWaRL3yX4do0foHO2vl2PkZPfoaY4EE387eiUts2xgICJZEQsrORp+dyk3
mWmJlMH9bo6IXc/g/7a8h90lrGfGK5fi/jBrLQmMifbeFTTkEE8VYPyDZN6xyuVWFm/o9wzlYsuK
VAlS2/hQGZ0Nf+9A7IBAtmJzJfjs6FLdGb5s06ZrhRwx4oOA87JMqPNfc2tRBK5K6M6gb9VpmOk5
PpikCrZNYhOhgVJMWoM8Om2ihVDpD+CDPISNcGhHMSItezc+7uzZK/C+7NeWy2d7fmI3qbW+k29A
8AbNZJNsyuib5k5UDCPrLEEjyDDthLBrJF6zwL5RoXjURp4oGxlsYtWtsqY8YMGWT9VLr2rrC3oL
3W59TivW+Nje6hIFcaMbwyAZNMWjfLWoz6zpX4ZPxkNVzghpBgOt46CpoINaDa7jvNdqPYoo6nVp
0mjSN/RwIzkQizlxUXZXVcgkhll3nxfYlFWK3MTVMoYTpPfAp3a9ellD/CUYhW9eVeEsrhajpShc
Foz/DPJZBU1gGfF3Jke4qoB83ays97FtjvQFmmZHxd+nxDvM4QAj1KIZQB6GubJoZ3itqyoKJoiF
ju1zN7oWW31V0h5sLpdbIMA3fS/LT2t0D7QsXVn7CpfmyLQEaTWrmGNYQl2Xi5iTkfCIFJwmVcM2
PTJEJ7AGUHZ9BF3h3Z2Walct5MLbRus+e80Eg+mNM3VHNG/xaVv8vCEB6UaGOi5yqvIAGKB2GqXQ
RDlzhAm/vusi+Vc8cOElyu70ufNRSIfcWfgRqQDp4BCUF3oEvqy4WEPSedO4Ep9x87TFU/sp59IS
x/cwYy002xk4D9LsxWBQC6KA4VPxKpmhGPC/87KCgWihucBScNwERy93tYwx90wc5/prNnuvhHuU
Zf9CPlZ7lN6lAciPfeCOvys1zwOHLpEVg06zcFYvaHCBmafrq0q0k7EK/TqMU1WSqAAiV9tCk+U/
mpkZzb9B/CGhoapKAo1uVFMqERD6Joue+0NFxZBQvTwWPASTNQMSwQvkFGFvwNx/6QxsLZI/3PtU
lorkK3M0hhEbdcQkcU+MaPSgVYOPqHzSdFkgUyquvfRDh8dV6uyDb+o55SG+EA2dFQINWtUUyaan
UaECoSUVp6yq9h68E9yF9AshVvZTfGfq/qZed/4jTWM39F7UEdubKqD6gQ9/623uF7r5WsYwqmmN
9VbD4Y9bxVea/tLdq2Qpu3GBwaOkSBHamBfsdXg+d9vwkGiei5aK+t4iK3XMz1MNGYdXL1jVGqCf
wvD/Eqo3iSOXc+XkbUKvAfH5DtpICGEEwS8+kav1zO0GjcxCVY68DSRfAqenQXBUDHsyOgcEiCRU
tVbtbrxjq3iQQpoKPUH+iHgVk1d86V8eP8BTCVsCPZdYYukanlcW+By6gncSeLBmyuBbZPOzJKvR
X/In9NZoN5zGS1O7DEez6+2lSGaxiCeT8r4Fswik91mOLIoxOtUlG+anX7k45Ufu9HPvPlhjFO9R
+X6kzU7SZRiwFdVYYDITNQ05GQJn3be/x90kyBScObuBllnPVQlgCbs29q41/sYhcQTsjzLl7g2e
YuYPpU8sUu+w0ljLL+p9Ib/do5Otce2WL4SGkS4iXVWumUig7uelMr+DsIYv6eYeJohC+J4mq4aT
j+QzZxPwpgsuAAnDp1duqkgVxJOUnMtL2QRBriQg+5VfciKuALvq0uG23DD3p4FiXWRoieT0Fchu
HDgPp+gb8iXGDQv8no2sWsHPGXKG0/uzYLmeVJU57+YvoRJadYGG10z/Lz8aVTMHyYPyAscXpjKk
0lKzBJUTGVSNCCgBWgVF1Vr8131aCz0qwaN8AlbfVnNqkvrqTKoVHTh49gpR3jTQXOiXBd8gu0p7
yGTr7pfNVtIRTs1b8fZvYer3tySbHh/fAUOWBDFafwyEY/SmpuG+KY8FzTQGPAho3zFNBZmLioDa
3R+HooNC7wH3jYTLAhXPGRtp24GDhx+DnOcLnxZFDSOE7TuHAsBcw2vO3ztCudzUEPhVUGkFeNsY
visinMY+1mhwiMrmnxakKN7EyL7VuA8BqXurXGjFFOQHJhbMfNlAI5IUzq+8kdpN/IlFusca/IKA
JyMQBHaz+lxi5B+skoJniNjm1K+xWA+24xpXWit5nL6o9CPgZWop0VR2yfEIxa3Fs6NNO2wI8kXH
vgMNS2WjQML0NKOpMqpseiNHSRVIRVHKN6ytdQvmIZIY+B1XEyWdWxV34MoIp6/Buu+rIZLoJ+wR
zQYa22QAqj7RmhwZx6T2xOIN1Y6Qszbt2zJobRlHdHgGSBLBUUAv3h7DMovP9Ap8nnFwu12AavHq
j3DB7DAEthlI+p8DI7lRPlrtYOJNIwqqcLDqZcOnwOTz7vRllFdbs47EbImYvDeUSARkD50Cc9I4
S5X9Ifj+5MCt8g3jd32BP8aK4FMEvzhmQKT3jTSJ6Qt08oANnpMFEDpfsmdDmyihUSRqJlCx2dw3
T25KqDVLm3mQzi+2G9TB5OuP/jCARQQP3zWdguCTFBeWxnWT7r8ieG2t6DoKkzq6uNh48houBf8I
ce2o5lh46MDyDlhxeqdBmDTeB2VzT6gDWcvbGd3WNI5dfkLSqiU0Ewpq+5+Kgdj3xR5sfQ+g2kqA
Oa5rBgm8pVU2rwuVrJLq0aBck/5A8Uh6XH8yrWR1V3x5qLYQ9IWl3GeiL+c0h5MNQt6mwIP1P8I3
FmJ84BSJT1o9Oi5/YsI1nIhM6x6hR5WPntSh65KO8WFtzcX7Z0tnI+sMyHVhCzUk8NFQ2oe/fnYT
dqxrvv/i8HsCfuqCPXHGmEVWVdy5nZOiOQFDfoGGyXbeaK2NESNQkySmozfr0XPr9kPA2yLYwmfB
IsYpfARK6py/VHcXlJb5q1oSHlE7Ry2qwMAl93MKhSsuGigZ/G1o3Ajs2Q6WXy6u/pxPSfjMhe3t
3M+mrzwqXLRYMmFsivuOGj66+zJsNGNugqoxwtlHm25c54YtAKRHAIMqGukIEm2/9+IHIe/tm1Tb
lgzhKWLgjDp2qjFdcVin0gWqb8jH5EoDnIFsBy3g8axW4JZ8GGpBerQoM7uR5tgE2VsxORD4As2k
1h08tPRtk6YhX+UD1kOr/HH1ji/AVZzHLMCf6S6osuq7GLJAgRg+4K4uOUBq3FT4mardh/uj48Bt
3Pw+czLYqYu8/43vHjPTDE4+vSEJhAO3jZg+UrusGR7RJ33t0OuNilVOWdDnLg+Hi7PG1PMooq9W
KkObDHGT4arI5Kvz+cYAnBURwrTyPFcu09n6zXIJMAYn/oILQ+eOBXh5QnC3PlwhdcKHGNUWQjnk
Z7DrzNUmvyAfbmAZE/DFHcXMkdmUSeKojBxyERUfPZnLMH2iUXIwx5aIsJIuHnM5l+rseP9eBslh
F/cAAwnqfsAqOo+WcCGrbGXa9kthhElsJNUKWtu3maxNed2kPIYD23LKmJ9pNt3Zo8XOzKyAA38a
TPe4gQw8FekOUJH8wdAx59V7UE/7y2Mudxa/SswMPN7mJh2brvElOVui1LzjjX6nkewIkKVAjEQd
TnoDFwG5v+qbqr/lfsjOmoszg2TgzSvksQ7qmVB6pmlT1NBuMN8Wqxm18swvOXSyaDDkfy+Qa5U/
jCQVSxTRLtCY4Ih/KNfQ+JRy/KtbDk7+z1cMpJGljVr+HMPZRsg1SWvPrSljwhSk9x2laSPN4M92
l2UtQBTYao6aOBeteyos4SlMk2EbrC4a2fe7DNDFsdpnt0k4ZiAcAnZxCCMYjTROJCGZM5qmbnZ2
GiJXt91HBg1FFFqyaZkT0AVkxqmKKj9WjyTDG6GoPi8q7kq0YOBBNYzicHYxMYOfpsek5bGmi3tT
0pnKBlLN2eybeaB9b96FFufLGimXyBz9ePyQcG+qnF1YlmDMunGY0X5AMgiE3unRakqw+U7vYCzA
osjF0bkm+QXs4JgBham+tFJn+0g7JVfjTm3lKCCMOel46Y2SfIZ0iGJ98KdsXgSZ7+goeIBDQWHg
l3XUUnYL3CwPIrCEitrcexjhiX4ObNplsRqpgWt/4kd+MM/NosX8TDnUbLrHXp8i3NZTM0SPg8m7
8EpWJUjzeBYFwfoQnV3Ftn3bTMwelep/GW3xxqp3sKpp4mw0Zc/L06zHjH1dqb8yGSPMlhpJqTna
9tuoDEu1PyKD+pQcrErzulBaMmaP7pHCw0OTaGX/JKdlmVpYRm37A/mD6YfHDf8M3z7wHwlCV8mV
Uc47W4949qEBgpzFSgaDfnX4c1hXJ63jQtNUavLp5P26qBm3+gkPpUVkHBFncOcpBIAF24tR7/Vn
PPyOVJgE9xX1EG1t7JZFJ7yXjdtZGm2/6pX9hB7QTw/qsALcN9H5V8MvxrKds0LBnqH6AqGyebu4
9+oGp0Tqyr2D630n7VVId1enjW58LnL9c946npj+zyJa3THA6TEqJPm6PdLz/WJ5a0/bWHk/Cb/v
9TI7qb558jgREO7czWssvWzSu02UbgNIG9ov3qIsLYhn8Qks1B4pTudm6d48eLHajx1SKfrq8EUm
0C1S2zzGzOvqDoc9K11kM755oHYPjGLsBkKXSBryRpYP7fMOkeI3ShmznrIM06qmBlUrROoxvIg2
W1rJC61KOneuiWqtIEkOHP3uBTXbRprQUAd+WUihY3VnCmT7Q9HDAYQtA8Lzy4yFdn0fEC2Kh3GE
INTDel6BQ0RsrcM8GhbVKdFX9qhjm2P69ladf/Ybq0hEItNMFnv7EcaTs+8qL+I8XNSSxvaxAgKr
/Twq/SMS7sdETW0kvg4FoseXg4UnnqqZJcrGnLyheUHez0LFVH1zNYfxHfQEY4YS5R8dUbUG/CBy
Bzeo6GgnT6rehWWhv9EMeKMuzF8kjAv5aUhGJ6AIYGGVdf9m1TQqjflQbi1g03HFsRICPnpioTwE
b3Ky8OH5IO9YYjJfCqHWVCBzr0Uq8fAhMEDRKFRuyH/olnz+7mokuD4XAU9PVLGSnI4Qk1xYsa8y
RMOpRlL6k+HelBb9YAX8UdzBURO+x6y39tsuQfIhyCrH2SGwUBNzXZqCQtfv1Fl6EeL7H2e4xoo5
EdAyrr3QlKQFT3QyswnRol4PSjncmlBVLUSmwnMkirhNgwtMCiLLN/U9qGy4rre79ZQyw6I7uN2G
Khx/8Pymkq4A4RqQ8Rwdb01pqQeLKEWDhFsgWdcSoOGwBmN1K99PuS4ckI88ptSiS065OBAj4IKO
gbH3bhBFNmDYaRy25P/BU+VLjE+1vT38/OACETFLnN7kgXqtCokNn2B09gfiofAB0mCvKD8Xr8Uh
34QoWp3M8doANGxpSs1JgK9UkOOnkwwJSZ0q3kQuLVBmdTA0gHVE6+XvZ48kxKbcBIpfGiaOI/Q8
AmMcWc1chxR5AjT5Ex8tfDLYgIxQgG7EiejaBxLGt25xNPPXrkO1iHDAzPr5uqtyJhzXZCED60L8
/Or5pR8KigC+m1g2yP0ldH3houX5X5BC7BhxxEFmMVsndyLkACHf9f4wMqoPC1B0FUUi92lg3yn0
w3G/MpWJXY8N8P1pPh41RpyPrJ1tmpkDvbPZ6EH2L2DHYnt/TFfImFuXNN0Y/H8NzoKeEY6fkvDn
ekYDUEaqHs5qyaXrEPbEwrVSh0EygdQOMLJ+QSbuMvtwp9QMazU0KEQouoMLjUQA2VHhNF3uV0Ba
Gu/HpdskZVY4z/pzxeuOLxpHWu6bVhbaf0JSCSBMM6iNPLJ6qnwnOzkDu11zQXJVXmKjC0O8RSas
jLO5Ggre5zfsi3eEe7e+ACEbR7i2ogvMz4hM8Ug/G/y0V7STzl2M2cYC68HYkRXG66JWSZIdpjkT
xRk4QydXE9F7PcT6RVcReq76oFvdLlA3FYAQhIof9q1wTK3GAP0IuTKqzFruCZKY0ZmG3oIiamC+
rDVIWBQ1SPcu1+nJGNxLbe5k4YvweBE3cv2II6FxO1u7oJ8rMWL1zRUClD9sbbmoJ39yrDq7l6Y1
YcGaS1JAzq5nHzx0tRiYGGSGPFEsSegW6o2O+tThLeIN/efNO6rIpRad0D8D1EY2vAZ+xf3dKz7I
6BOfw4eV5udZYyDuJdsuKB9dK/fmNGNQvnWs69uWk7BR/Vp4y+hbE+KCoTjYXyWdIjcQnEMQF+12
yGGU4TJSv9UL4z8a7kSqrq1J/WJGVhZJxJmqEb0rDD1LanO13JDgBKgfRFVLu6o7CMctFdOCggmR
/Z24BeAABekeN6Czr2dHcj3j7fqGWwuGnfa3n+SPtdzjvhDLT4bjY0JCFHkpe7mMgMVZHoKNbvki
yGljPBY0XrV3eXPA/cj0u/F1iT5H28Y9SqKYH/3TcnOcAi5RGdZ0gnKXTPLbGyJVRxdiEIS21wP9
4IeRuXyUHl+Mv1iM+7hPNzoLpXI0nmLEBBS/KQ5mdyDAB3V9lOi+8Y914ioZjVGBVhVwlSuHUNCQ
PRKASV80xP2E1YHIQX/nf9l+2f4cywO/GLIu27gBXhOdi7Cc7uFMZ2gd3SZTUdCXibdSWNg5lCNm
8H+qJ44EzStknIj8JEKw/tsxYEEe0yAkyr6mFOrCH73rYgFnGzLHHw+JhUF+TdFxXCiHTlP+FQtW
+hEbHcQOaiI55HQS1QzBYO2E3pdDnO5/o70aFUm2pAXuUQku8NHUtXH3mzm89q0Qxmiv/XrveYET
deh+N80BTnGDh6IC7C5mv/TU/gF7hZ1q/PBW+U1VCdTWrUCnmsdf68dUM6n7lQyMrB89J2QwN6P6
VFU8jdFUbIkDWsblT0r3tm3rWZM/wwX7/AY/o+3Yu9OwSHTFju/dmZpOOEoOj+cRj2rsUhQK1ST+
pRKnCtW+m6DWE/FYYD02bFLn3dA9Ay/53g29qhvfUN9p5JzdH09vhdRPDCQ+kcwogDRfXy5LuO37
59k2rerLib+safOvn+ky2TSctnxp+oFdFJUEocfaZ5/T8RFx8jgr4cxFdqwky5O7vcuDS4DxDhzg
b5NedojHxC1iR3cHAkjGbgEMykucM74wwRfLNicWaRJpxi4QL8bkqilrriTQb9b+aJaLuYB57xpG
NOj3mAD7aOeFYQICz5G7OqvCvKgfQeHnhKF5NUluhGAkk78zkMta1Jep4wyg1qn+O/ahWhukIdIr
5vRHczpwzGk2bdmSkpRNorB+2pu62GCq+h0EsRlNLXlzfxOZY/QKSbffJ3tbmelwrCjLEYFdT60r
GlaUMMo/RC77xh/WmOUBhuhSXxroG83v9oBdGuUrXnLt08VIo8st8NoFY4EvkN2Le30psHy4upKs
ONdvQHjSQrR2YKEQfh8z/ij1Jh1E0U38iUKw+795eT8JxVduaZ0B3WodktRkDDA7Bc7L3CJv14qk
eJLoczdU3TF3EX01T/7EzLRuAksshF9znF35mR17PxtbIinxp7XP8mLgYxiPB+YluUD7m6i4aR2H
xHePHDslkSLKZwYO5qmH874ou5ffsyzR/UdJLsANMRFHNPiIdpTvppl1uGEefazPeL46QR9xBSUH
UkWRz4D5qnhOfVvcZuDEPGLYKZbpqsf6H7Hu0z07dNoF7Rgf5O3vTiSkwiixefiZRDCLVP8B/4Oc
9jPaMaOVmbIg05fPBRDJx49sCDvS3aLADm3gB5R+bxfoflvsoXVrdiqHsm9RtALxX6/6WzAORm3r
JkNCZAnOCqVD8iLVdLO4ndL7fFAdKglrZMBcqiWId5n7pRw1NZ1Bgv6DObkwIWk9CEqYjJQLBW1g
tky9fIE3iXjYlkdmBc2xzwDCm2ytamVx/FPtaHqZcibvcOIUPt5eJQf7arWtuGnkSC5MKZ7LotFk
cGrRtxcC8X2waNS9YUJwTN65c0/qzXJEaMRHm21IROK47b3+ryKhLz1ZiRiEOCUl9GnFeoRvuPEN
FLaCnvrF5CJ12yYffes4ts45E8Hr15oMpCVcJyfHnOvle8OuFKvIhaT3u+o+N2VrSBV4nm4jS81o
K6NlbEuT1hV4UbPgoZYRbCX1eXRGFYF+aV+umqQr2KzORc3cyoHA4ewUJwKunfU1fqPPpgKFwZob
3BQPbR3KtzX/PWv+P6Scp7TAsi/jrBgARKHXz2+RWiZDmQCTpMAUBPUWOsQcqg0qjVomgmeYfhPJ
RcjK/qIuIdaXssROklI+SnXoBxhGSMVtRA0G4MpkZaO4u1QHLmYLptK8eSfjPEUQnnhNK/13RHzc
HsFhOO2KvbFjh32yAUODtbb05dUgoiLzkprHR8vNFDAQrI9QfcH1n1KQLjybQB0UKd5Xxzdf5hi2
mhVJ7ufNHCvyjTI8P1ldptpVPInfzZZfb/5Cq2pw2Q82c0g0Al68y3y1QOUb87IN+Xo5EEllKngC
X4lPCczmxZMaVUtb7soHEhRrANV6G2Dux1m0flnMVr7pyQdbmU+FuRLRe/Ma+CVu5z77zmKYqROV
YzQW9zOvBkvK7k7r0ZP1QVMG2mV6Zw06rs3Wk6zdxJQWnnj3iwygCQxvSw2Iu3xbj+1iq5VkVhg1
hy+RWIKRD15JTDAiOfKckSpB7wghOTCxOoW+OzjMuEsd2UdplUFOKV1C2rxbb7IYIkp7sQAZ88h2
yUoazWJ5J6bW7+wF4eQVpOCOKwBesOV3IvGfmnjDEv9uO9Ou4znPpVaTh2roHAdf0Aziw/NlVLiA
Z3I1gy31B1rkfhLiI/ZLyb/ZZtrdwRLYEoCRLSp03z/s5OTosG2Y+l28wKYbAGjg2ebS4ydJ32Nt
RlkVy6vJwmHarqliDqaTMlbh1wu0J/c+eQpYjfFiZtTkoKNok9W/Gf0+PXbCUF5DB6kamRX6jex/
9u6HVaPR0OtmPSLk15wlpwrodm0aL8CIx0oix/bP7Bfrzk1CTXEQzYmuX4cbqfQ4rL7w45TNBwnC
ahSbN0kSV6ZgPpZy9B0eW3rqsK3JmIamAWSDnbdVIOT3ENFRfFFNCrGq1yHBlQJWF7Hw5uXRfDqN
Xw2GN8lzlMOdXvWMb8qVoQICfbD+m+SSBRNE2NWfcaJj3QuuH51vS37lJp2Q6CO0GNRBVdhl1/+v
t5uDExrO38rpoCwslwJx6ouTaja8dBs7V3wgf1l5JkcYJ+jpHx7WXu0z5VklwDIfE8MFEHQc5KHW
I+MpmGdsmGE17iA98k9S9eI+9uIoR5DGRHEdBgZrqsYwvwnSM19ETIE+4SBBEydMfqYc7OKYh1i4
I+bxyt2BqQHRoBrqMlpcQoXL+0wdH3KCf9AvCYWSEti7Jr3EAxEsIDEeQjHn++DaXjfXqA0Kl7cz
Diy9AMdzYAlbiiZXLXTuJShcGAbc0vxhvUOF6ipqnoB8ZTbSW3NH0M4FVi3NG/keuEKGqfYU96zy
luJDCBvehALUyOS3uloeqc2GGIHhJagizd2pf3XmmrIfuIxaInci/4jXMkupfHYSSPrZR0H3ZtA6
LDkZS45FUoPpysuAWtRsZ8hQ7nO74OZv3hfjWjtTcP10DOqJNlGEfzrqDDXOpSydmOf63k5F03IL
2oSv1yOXRRdJIulzXVigZouwGCxAtLKS+giXmkS4Qr96aSB6jT63C/yvvOPj1n7jy+DbBbi8rL7y
x7KGn4erwP3fTKK/xbhAJXabSWBrb8y+rq5h4lRnoLW8ldDwkuTcYHuOnZ7iCfJiv7GjQmZwGv+1
LyHcC5+udhsOKE9KynWuivjWADus1LJ/6gGzuUsIUPa1+hVC4Vy49Dv12ITIhyUi0Q68n9VYTDTY
YWOBLmfSkpp+OSOpk/UAHPy0VtHRGFusesx49ch2CojBvPQDYzc15T8Jw8eZ8w8dYIXOisxB1XN9
HauEqFhsdTrmJ2PG1hhDyDl5dr+ZcckFxLGcY3+rdegknD+5uCsTCkwtfjqKDPEqCvuycfZHqdRp
cUSs4g6SY8przvcsYi52vZu+bCDZ+ZoS277b4x6oO10qds3VPV3umLNdfXZvkFT9MkZ7qKMulDk1
rS4q7JBoXwWGJO6LOM2vWDjGWVhU72xTusHjcO8RMFnd/6bJiGnK3BPCVGwzF2YxEK4ROXUgtGy/
1PFtXzy7e4fXrrno4ef0VisYy1j1YLOPOD41AkJv75/cFUxfCTrIWz5Xqx/utn74io0vFWt4G43x
836tGOLL76BSJo9qSzFiWL8YqDMC5VkWN18HXp2UXl48QEXN5ut9xE29qY8PhUV5gnCthaRALopU
OQR9s6CP5jQ93Xx569EUxINxHaRfM3mLWJUst699O9hdxVxlpmEV7xre9FKBXBwRTuhUPQanyRpn
xGZqn8ZtgzungVYUdRE0vCaKU8JSf3v4zBNS3yOyilOKGS9YYI/CDO7D/3lNCADG1Oq41qP8kH7+
qlfF+i3lMzrLW7wv2a+4jFqx98TRv1yAlaZMjNdy/iMG0UMZwTE1bGvqq1JCfcNm+9hiGA/88K9/
4yCh+/K3b5I3aNy29EENFJ4kw0hUslNtCEdhmMuiwjflATITSFtyus0IYSQ0Bz3SSP7rYZhnVAQ2
l9Ee6OE6fC8IvukEt5hjBnHZfkak9bnwmm192P0daixOxWN1TeC0kESi03E9Q1AYfB30+rFvVjAQ
rRWPEfH1OX2YlVgFQbBqiWByS8rRQt2/DL5+vAx4X7VW3BS9DhAxi87Celnii/YdW/QVaoI8WRjh
e3QK5mos+Te0mGImy/eJBsa2KtwXfgz5Pf1ZYIXq8t025pNuzQbiq3+iqLhIBZaQ2HGBWWUTYmk8
/CVBIyFY+RksvqxteGoKabeGZCtha7VCSywSIBDLQeiO8jA+jLbAHeLwrbbrPPNtFd87DRP/dqD7
tB9urPXvn8sU9jEooqIuMbRLrM4kX/+ljk0sHomw0ZJzIsXGeOPSYOUhmJUkRrmUeex33bd3Oy1L
226R7IrYWUyHZhRHMAfbre6/yXhj5fEIHD3WsHhm18tnf59MD9hZhRUhkp9sbRU3M5Q+8sF9kCEE
w782yOpoiM272LJQgV+LWzt/a+Xvkn1OLHUDfRMjohdVQiPQyh1yow7kycseuDLvM04KX8Wyp3NR
LQ28vTn44b1MYtZUTHEn3HSmpMbtv79ft2f6wkeXQ0C+mF/ts656+MmeyGA81OXwMziwUn+lmeB9
Q6tG09TXOP3an4cW08Z/LLrymvBrzICy+4iQJwWTVDz8P/Tf6hpi7DbKbHX6F/NsOQX1jK8yGEoB
ja39e2LjwFNWuPl4/De8Z0LA2PQ4XC++u75gGWyPC4j6n2eqM+cljHIOYJQzL0fDAhK+MK76MHGO
n8F7DBLTkDubfvDobwLGXkcbhNqqhz/9USWyna/09S3dFX1CfSicmQENyJQLMbC6SOGso4vAbAnP
LM4/psGaV84Aab6ZCDZNXsy7CDx3OTaC8Eq6Oh+crXzHTjN0rfyJeQW/tjlz64uxxkCGXyACTqAh
UdZ6NJsjPPSUQGxEULOfTrOriRbbYJgkwmgQ80uWUKFwizgeTIMx3oBWvGpr3m511e/rx+1orAdi
OWy47gp0PaywJjKXLvoFHuxDIOvITmRWVy81rYCbBNRAgYScQ5ntMOmV8Bf4qye6oqGk2FYezJWD
HXgN5Ydu6aRunNDCwu0GvFMLEeOV2n7IT/S9omjktPginarD7UkAPOcwxknCpB6JgTDbyj9Id4fy
nFDq7P6/CKTiFa8ZAedqiaozEweD4ikRP7BU0Fqa0rbgT5tDLS6f7Cv2lSWImqOjWsJTThRA9eNY
tchku5x26r4Nhf2fpWONh1ElVIHRT0akiJpM+FfrFYD11qWQbmRh1KksB+rNqwZWPj8MlELlCZeU
4co4fD4efN/n7eLs8fioxuRfqagd4MgK1eYlkAWy/Gu6GA1kqswqZipWYZ84XyVuO1HTein0cTJS
ERPGDEBTa5GnSlY/YXCAMA9CGqDCj5kGmDYKSo8WhwUWu+OwSTgveRmkj9xb7xtmLA8rlkzp1pod
tuAMa4D42ru+rYzd1JwvirlIQ83bRpnWH6ZripZrj8q/RswLw5g+SQ/X8O07VCPEiFn+H9q5W8Yf
Ai+ImQlNDDaXB0Y6FrNKKa6AXLvOQlY6fv+j/g5x9nUQHRyqUzNgPICrlPuyHEjJIOuisTU8OqAp
1mMVNOzRFYJTffYFXcwhR5ujXyqh8EJMhjkot9YgEr4UHE3mO7Ee/u98DmbimFj7LqEJU3C2bjEH
oB81ZRnYtmiB5px/BUxspxolUs7PAvBAyjastFAuEKhkdc97Vir1XsO6LVt+a5hc2q0eqmPcH018
ckU9LxYhXNenTp2ESbXwQrwUFOPIkLs+wXziT9hlwYvk7TXnePeCSZ+DAu4qMvWmWracjPcXFhaK
0B+SK/S1SPeD13GAVHlfhP3Vxj3dy1fjxwLH9Mo/eWc89lS02lygePU7B/cXDEPsFtyTEGp3SpT6
9RjnvICczNvtKKdA7zikRzEHH27qH2LcTarFVf/EbHGFnebjL3hW/0MQPYL+mjcTHgzEBiBVXBa1
ecspfIxQ7Rgz+ZhQTZzE0Ujj87wu+Q0kXzTSmhMjcqkg593GpLTTDKdic8NwbGbEGyx2lmK3Yvrh
Yhq5or4ob2/2Ec7oIf2rJdwVR3S283M8orcjSK23sBgUBMxySrgZyDxSUKmfyrCJc+2x7XQDAd6S
GxEkkZ6qakNYdzgLbDuGZOjvvVQnQxCS1J4dO4SCVu3S0PViOJ/+cV6E9naCfg8732b7HfrghBxg
kZThYvzHCf7/od7HPeuYnvwmmCjc+Jp1p2fuRq6Fuveka94LOnMwjVoXA8U8P9uTyRmYtTcICaJq
MiPHimzHRQpQE+QoSpwzHA4R52mZ9Fhc+qpPI6fNCcVB6ZXcsy8KFhfjyV9L3ky5kuCad+qFJSsp
XXJKsz/5VI7ds70+9Tp2jzqCI60gNtaLJTa7o7AVtmIT3KUoo99wM9cuNhzA2U60JlIZnVYKQOHn
XW5LFY/vNmF/Sy9qrxzBWP48qcNGSCDgs60cir1QiQ/haNdJTHfPqqcT4U0umqSA+kpIL1ITZ7lc
iQJBaCUX/agq/odiMoP5qBeYnuJo/ijBdLDvcd3ijHliqr8RrVJkOaW+InPXmrfvsoA/2ays/n8Z
UlB3j6J3ETFRrL1KUacmu/eN3Aapqi1Zn0/7Fd+fmv1nJ2SecmakK3EcR6JD9kiETi/QUXDRBNvW
9+y0bLAN+ZCjy3fWweUUE4Ek+c9iJxZ4IngwSRHtnwmBSOCdyTJrfDKIAy58hlXdijEzA8tLVX4N
DUU50CU50nKRCHazxU18oyuq4pyJRxSVPFoVeJO92+Y+8O5uhCHh9kKlqJb6K1Eohq75NTL8FrxY
kOgresfS71jaQUq4R+FA57XsXOy75h4D3eF2n3opE+4pDFFRzpaYnjE5bRWGXaVEwxGyVdgLG78l
UCOLIf/aHoYbtRdvLnDQEP+j86PIkraGhm6z5dMfV0runCya3NiGi+XhCt8XEDYHADpNiS6nJCD6
tsU8vsxqfpc+MviXXR2iiytlxwH1wuaL2k3LG9gkdtpbDDhPwel+RpJj4yfqQe/AQ95l5pA2R4oA
0Ag5F9NxVpDuWCnVgVpiSbrrYQ7C+rav9xjGTVBTBryJKMdsgdeKccuN+JWrmU+UUNUwfr2k6z0d
W8XPQR6iUnf6NwiQ3bPs1QJIH3HnG297qP4nQOzpNSJEWlA0rbxwNynPMbrQGdiG+jtQ6B5bcodu
mG+43LxvH3m6Cc1tQ003nbRVn3vqAfBrr5bsJkO8W6x5hME/7yunipZMSokge3TcQHLQp8aEw2+1
MGHimoRhWf1XJaWraztNuLgObj/suUsPn6reV8O6JCryXrkVUInQc0fllWQYVC8ARGzUFo3zPSP+
aBtQSuGJFHwkWfjShuI7WAIHZjZqY3hvZPRL0YnievHBpU2kwauJ7J6S65oPm87okebDfGPcjPiP
0bQD9HUg275Nj8XHhKGPMwHUmGRxJuBkqkr1gz68c+KWZvrgUvoGAHRcqfG0RcNw43ibt7zHPklI
ikgFeoYQIK0X2s2queBrnpcMZwAaeLoJPhNse+Yr+B9b4Kok1Lmiemwc6Rrkr0R9yAoKnuSEjQD1
ssyyvICmYeSJJYVkN+g5X4bt9dySj6Xz49tApjvZnXuBwNOUbEctP0wuzod9qcZj6EK7RYtBnb65
q2bJpTKNPlrA3/k50BgV1IR17UKgwVZ9PyvvJks7QROHpuPWERWy6ohoK5ZnPAQsFkteW5mv24HT
vn6W0y+9cB9G0I5qLk59kOGhW3y3n+jWt/K4BPG+pxGkEAGZDcWo/CESBmIOlsg7ozYo/I7rPB12
Adc16MIbbPCsOwPgYE5j2NuXOmwispRNSJXWo9y3DMFfPZEcVawSaPr0XHeds8hQGvxh2ewZQou6
Ebo31Z8lF3zHPC+JlT1vtnvG4pGM/KrjUqSpnFacZsjI01k8MATcHx1nvDSlBMGQ3PBUyxcf+d9r
CZU9VBoFBCCd56/wixmc8mv8oL1EbZH05GqEJ8gqpredBj/9wMobiDI/8PE9KyNv/yWLKhATPJmA
XJ4WUI00ptM6L+acD+Rvt9LOm8yGfCiEOtZq8793H/wP4q+aW3zXNtCm1fCYaV2l3Q/gE8qZYQGg
793d+4UfalCtb4YJHN2veIjXF9iFMyG/2L4/Uzv0uoHCK4OIn7sYYT1GYhYdwf8YatSYDLQpvajN
D+feaTiNbnz4bMR5E46/d/vD5jny4A60ofPW6bValvVfPqVugD7EyxM2+7b9gOVhi6vriNTFwyDd
0t50GxFMhQtfMj0iQrMhsK5ss8Pj7b8dmleEbMF4I34FN24c9bJhNdra0zpinFHPiOY+hwJ6NF0h
NLE224vKuzLPxGflQYFWr/I9If563wYXmSxe70Qajl7Rqv5/ZX49anAopR9iQcUqNknIh9+DckMt
U7j9cTO8V0w05UDPYdkSVgQOIU8Dsx9yaPx5lRZ46/ayJ24czNGLcT0ZqP6MOdMliiil4x6i29/Q
OwNjuyeYoH5T6/PoYY+MpqUZIr0dmx4o4XkGv8MfogiIF1x7fYlB3mTvPd69x/JbGmJ/kpXv6nJY
jv7l9ZlWFz2silVw6mOq2WhF4izOdBXWDil/DEE7fbJxT9phB8bu90S4BOFtxVFTg5zbz3MV8MQb
itOkOToLWFXmTHk5oJimwwzGvB0VxIO1uc1QoIFdaaLyBfPRhKvStlgLog1gF2qgt/IZ/1uPgYph
ZKnO+x5c/IgQcNAmHM9K5YmCVYA0XpOIq+qZQjIY4H0AQBOScN/mlAZl47eu00qEt0vnRPbhz4pr
QgB6kal6y3hU+uAmNn0qsv8PjThm3R6oRbl3tWFFcldFt+nA4fIkQ+PjZfmCuaSA7AfPDcwwy+px
hYRRF5pOe342Ot4FLDjjljfg4s1T6iQUOcgJK8j5VKiUtiO7uDY3g8e02KsDNxj1mQ32tauSYmh2
qYQUoAaihvhcivkU+OkC23B5GNmJ0I2z712mZ0ueXXPW8SFJMjy39JA9Irw0vhx/JlmlcSMCUUeU
Yc+0jymax/M4Bgy7ffL4IC9hiPGEX7rf0XW4NGasWbB0vo6Hpm9RpXZtlU83ki7K4r2gnCXEwDqy
AR0xrfYaPHSNPhQX0nILeeWPoycSCWCBFYkC9UHm6iGHs9gPlKNOTvZWzvHDJUYw7UXEt5aQkzkp
O0a2mSRuOFqKZBMBB8MOCDdqsSBkhGNU/LkX2FdPU8/cf2Y9B+81wQw5qoWRrnVhbnbO/KzaOV2V
+nEaoDA3HZKqLvVdg9MTsR1wGxCKciNsHWXQHi4YTAstEbtO3nt0895fvAropPe8FuD4EyVOg4Kb
yFjQeTjussRAAfBL2OXNn/2ygPkrkiaiDIgk6Ibm1oeO8jcLMt/ZM7cYUmljbc9c1clarFhRByZe
HSmhtwWWtFmjzaMfH7Qy/uJ/WGuN1RS+eRWARwmBMkIRnf7PbLQUdoWqFhUB5w2QTMazXu3O+okh
HDBPTOkZ8RxyiagOrRkj+GNx99FCnRBj5cILwq4EkfMTI1KjX5Om+t/CJOXqSDFBL0r/PgPuYCkK
PC5KWH84wR53bfGQCa/HYI4u/629vz+92aYt2sLdLryNUS3vOpxHbPeIquH62yJpRCa2YLD9WxTM
exeZYJQaPCmh8InODhQ6eAs0mHbPcXhtdXx+i+Dmn57xCRNTY7kYurtnBrB0Yf4+IB9cvKJc/t5J
P+KXSBycQDE+os9vinLZKzOBDJ9bXtPhCNMK1Qi05Jp6FPeAmKnrZeLEQ1Xx7+TRvFgE14U7oWWN
tWKIRMhlWfmmnkogTWuwszd5EDnE/7f9eLtkvX2vb73oEwmxb9tOHoyrLyBE7tu3nv8VBRnRz65m
GeNIzL9FCU7fpCi7CzEuEr2Hbg1ihMBCslYtLVE1HqSzRZvq4Ttsg1Kb4XwQ5PdSbHF1Fmf+wYav
QA2ZlDN7ZyvWVT4Badhl03j9ZIpmzM9OZ7JPBVVzz/izsPqwAG5LvMQpX9MPv47AnKPKzzfYL+xc
r3LtbG61mrSSl807CXmSZHwTkDeCFRQkvmIx+6O6SjeLJ5JKdgO1MggDp5qsbqD2zkTmu+j3D3XL
cDkFV/gUczbsh4dFyLuJHK2N/F/lZsQzQjaJgMVPfmrsvA8Avc8DjZEVWFBTWsRk9GUmYAug0iug
l6xMyaknR/XG3WTbuY5aAXGHEiWO78N7Y2u1yU1dtS+8eB2w8h7d7eP/w5nnT2Y8ZXjCv55wIcRX
btgVJTqppIb43uM66iARjDeslfIznFq0KBSkXR6TQYP0RZj8Y3vA0knanSQmLEwL6d1xBPaXXB6+
DyQaApSnZ2T47nt3UHWY/JaLRZ8uLPkeAlFyX4wn+fSoK03vhqFfHiIjriGJypeOT6+OJ9WwnGUy
6q6dai5TZqw8xBjoiiYLv/N80+11TFwOq7U19nNCUsPk7irmLq5irD86vrmAFADkB49GT5dcxmVp
Bfp0prrd9jE/uSEO+dvUxUSuPk9hCUDN4+LNM/BefBaV8ktV+mzUi6pyOwm1hfRo6BFWOyjEahsA
w/4ltQ1M7FWFTSk7ZDrf2XlOB9/6sOzVo4d5/zqMQCjkKN2Rub641hQDDaVzCzW+6TH1gkzSFIZD
BydWxCpcYUG/FHYWD4Ko9NCgYFnA3fGljnyu85gYop6UYzEcDqvm0yE4XnK4A4ScqJBFIlHOhJVH
ICM/J1c1tiWAGZ8cMQ7lcuMp8Xp/AIXgBBhwztgGXJ2N75xXBlbEtFoUdXzWWZTB/W/NBgz8fpHI
tI35z1xH0HFoFnXNVLBIIsiWAgyjB4UDvc9EvdYMpDgucwIJS3Tjrcqau7ha0W4kXXYh2cHV5gzN
XBQMIzFEzeujAWnjg5ApbclveZglIN7n984fZP6aeJVXsOVuiNQvjcuh47R2KTxy9HV7yr4Aj3XR
ZIYfPZ+5LJocmcbAksYazI92MM25/A1AcDkhzoCYoeWbsyjtHA8eKCWnGggMkN4imDcHElFcJa0i
hXHpafBm6dZkKBCjOu6Q1b5Ik0Dbvz+dc+pcXp6zgLxjzu8DXE0McqFfB6h+kvcfRlzUBECapC9d
d12jb9Pect/jnI4ylRNGFnTrKsxV5MhI3SKqDpFqki0cc2Bs8wFRPJamMorXRtFf81oaODgjSZlf
SuriQ57E57HU/WVAb9au99csjzG7gUzCYctzu6qUAFKvmHCbG1pSi7JZenaRBEPPCM2246jnSRoW
rw5rP4/YcFuRgD3RSXs8pOGeMZfaSQG63XYC/ejsnvW2+gipKyHrIEqWjYLQoz+ltvJmPRpQL+TY
T0B7fvz91mXYuyr/sz/NQYEr4n4B+Z82IyKkNK3i2ksJ+Mj2inS1GVmkqsq+58lk6iK8AAdBs9eb
yEQk+GHs0HYN7EYSVkA/PdoB7z98P+ubbHm/anH/aiIk3grK9aZkyFejtbnYc9ALFvnNJ3QAq6by
uY2TS+Rj1MyIoAPeVHq8jFNtQr2hHqSDJ/gytrExSOSUGymkjOXM5dqkr3PP4avQOJ9i9+zRHsux
5eO3LsxjCyR4Y7R96ebNh/chBRMvTxJuHSvwV9WmNh4UMSg0IDtJMM2SVlZ+nB+SG0eJonaslnnh
qeRnQnS191M+U/vs9fkZLlFWw98S8d3Z76OVVascQBw168c9fF/ZcF9H12MjrkJzRu6r/AOPfM1l
q9JEB5gdXpVv6MjZSIxOPmsq8yJNSmB3+uUZK1MTNKcwnTo/LYJ3qSaeZyhnvq4VvV/mn+mIracQ
HFc1ewyIZcKlTwg8zbDbWNjoVdJrVDOOlBVwUlT/i820DMKhsCc0hoGfB5AKl5nR3Iq0xnUQwtNQ
Ls0Es2N+ScrBPg1eXG4wndX1SF2ckPvnFenkd5yVdaIy0hO+qmVwoJU3ebQLrxMlF4AS2gS3j8uU
SlUOCqr9+x6r1sEdIaQiF+frU1zPo9x+kBSG4hEigtoWnfxvwGK8mEFnM1b90hkzDI0EPtZVU14z
HDtDbHp3NX/ZekIaHH9I3bCPJTZR8o8QuCn8LPHxVMVnW0m6x4ZT+7bjM/7McFYHO95p2P3V7PVZ
EMZ09ci9Q9Rl94lmVJKym+P4MvcSO9Ma0NB0eUfm+NB3lqc/Mwth2hMqPkVtxqOq1DWnq/Zw8But
VAYfsVP8y0/iTIkQY6sGkPxv3byxskQbC5S4KURqoAI90OpFxxk+VdafFkVV7nLK5e07s4O2PFzu
uEpcyOE4+nSdUHmRkMwqqMfGeb0vUunYUtVEf8oI5aH89xd4MtlSxSEVaq34aZttlwoMN9PlKYmV
QUH+jpvIXDpwOuNYrIm367cQQE7Gp5jZHkZBWLM9aJyMxaAdnxfIfdBNrNj0BoggrF255MObg9KJ
eRM8T53lVTgOxeCXd+mZm3xbQ5GK1Cg0HJEYTuJOfafJwW+GXQfDQzE0SQ0VMWwr7dlginMUZNmh
Vexa6fZQ33ePZ878GvShWR4I+PdU/9PwGrkOC22rbtyf1G5Q5+/mfPY7BKEPbbs7CStp2j7J+00j
sTfgjqWEcrifc6zdhQx/BIW6XYJAYf+lt4JNKX14ll5tbgkbTzQezZDrEgS0paSNj6/B0T8UdVie
llWaXM1xS1OqpOovC8RfSe0FQtBZr5fle2L6SPV0u5xU6Z9DRV2nfHEkZvCLUypvt8gujy3YvWeh
xxoPqAs6djEnBKyWjqcSbeUggzYFXelrRaHuvrBVvY3dxr37Wf5fvkO00PRcyFYkfPfA1Erkbl+Q
Y7OMcfE5tbTOR4CdpWmtbQ/0C/+CMFPw4gVkX+zsfdJ8yNord9xtr3AmGjIqSkG/kMTiqjfAYVLA
ygezyM1vXUtkJoW39UNCMRZn98ZJ2wCIRWtbNFu4ao6dOwE+hP8TyiiOBOY6dEYA3vAMqBgydM3I
BxTFf9SdjnWMh686PXn77aN2fwVCfi0X6hhoM3RvPyCpkN1EtH4HMNUKJUz8jzJOHwmzB7Dd1APY
A5VO6YZ9VkS2wvvBuOBzLcEXy1UtQCZzD9vPXpGYDFuvzsQPAlz9Kcsd3cwBGreHFTZPOzg14rSJ
YBYhKmUE3iHTOpEOBNdLIWPSCtDwRRnc/Zq25AfkagASrELHnSq8+6R7obtuayJTyeZFBpNNtydq
WfzJdJySMBr9oRGM/0J/2A3O6khHv+tt8OcQNTSR4NsqkjLgPBSJiN0z1MNq6ncrYONPZnUWXxdz
No/y3PK22Ydol9/i3Vu3k55l1cER/OCwUVihAjJakXdGu+JM3fvlDQeeQD5gzWzQ8h3y8VFLbY5l
vJc0tEjFrA7u1MGzKchjxby4W6kt1VWoV3X9fPrS3OpOGOpjdIQV3hXW3r72GA5sorboY3bAKLr3
muv3yXuxBoUilPB+sXvnliCWA5ov15MRQ/qX08udPVW19z/6zjD8OVnvRE2Vd6eE1F7DrTU3Y16l
qad/yd+at99gu4U84HRiWWTs69907Gi+GL17GdnuNs+OMUDBUz6F3COv+Wz6GT+5IY4NEPr6qFwO
3bI8Meqg7px+oZtzJwEBGCvuaHWs+/bN4+imgcU4rQqPDzyzf2ynOLMli7bpHrBk/hde7l7Rp+HJ
XuBA7itIWBbWslEsKVBrVUInOJPXJ8ImlYVtRMSgy5/bHqfH1mh0X1aKp99KBw2GFDcsX9aZ5ItH
qkkmTpCXRJ3VfPqWSFGyOa6vCv1K9G/dR+hQ7cM6yoLGQ3camFwWwKKxPL+vyiL7fDSnxKiAjIzA
LpDKYtN+VSbSKLxDOSev8Z06WQ7ZplogBw1K5XqgRxZJ+wMjeg7ZHLo9r8NGtk6FOIhwBh+xf1OS
ImxpOjcOGd8hXbEYP6rkfEDc236zhL5FlVHSHEsZSqD+eS/SsEBFoIjlLZay38ob1q9Ryxf8TUrQ
RPgA2rJzajt2JwpwgjSzWVCsyD+lc4fqdGlmJBsLnR9nh5oWvKrPJfOj+p4CfcdDERl6TunKAUva
O6oADjF8O5PPNG3KQHlOVc4JZ28U+hB9FnwgxNz4h/BnL9XGPyCH7Tsw77XF4C3e0HYAhuxzQkJc
zRJPkBPuKdgCoHMX6eJ24eZQxHfoAQy6ERah8G8h+DzezKVK3G2MmruIBxVTlvXjEWzoTPo4sN/9
zGXE9ZvhFIlur5QoXYGlAilBeXOVKH89nHt7jM6l3shBaKgSZDgOAYl5Ie1ADNJrdOcfiXY9yjs7
8UTCwjji2lQSadNte8azQWJAGe3LS8gwJVlPnnXGHeyYoUmti8kSAIQPG9zZ+0Y/RP2A5U3WyWT+
63XBzrp3+5g0aeX/U5kmNrsC+h1YZ1+mSvvl6holKHilPjQPako3luI40fTI69zRgSBQ3QPGTfPm
GrwIx0XU7WEzpt8797mZHXC9GQKMt6ENmE+Hs3OiGSBGbwnH2IY7d4JuT8vtF5glj9NGDZ0Sw4Bk
jMQ2D+gJuof4kCfKRWs5C4Nb40JCCKQ3CRn5DO64BPGch+JyjBKzXqrrEOSkoVG5ew1XE3ZGS2Og
q55OUZOjEefMjV7iiL7wGd1HB5zGRTd8LM+7CmrNBs8eX6OaKy8A1nh3a+ovy9nlc5ncUJnvLnyb
29/ju67kTOotx3oD2CkLEGvXoq1B9vltJflHtTftnBeTxUNSmjgyCbSGjIEzq7wcPBpl6Uh/vCiq
+LHVdI0VLUhaAJ6qfpeMDtRXwtRl2XSb4xZYPbCQkW6UeJhm7FoGuK4cLeUL8DJvrwYD1XLflFpt
+Hoi7eO+0TVjimqiP/ZkquCcm43oL1oz6EyhbQhPoKpxp6VslbKUTAECTg2Td7P+8hf1twPdS2Eb
7G0lZhk3rMZsUbK69uFPyOR6gFMwyy6idSIvs3rBugw/fyr3nvN+Pw1ZrpOwYUZRoRnViAi0spCy
+10A0sr77KD9ZapmWQO54gOFPNSahItVC3pZO2yKsKIdQa2IHUWfTNf5TTDWy7H7HWolESudrsfl
fVqq/q6NRs22qxt8Lb0TzckkuSww2wI69aOTKQIfD/+wZwr5vq4dzkc95AL4/PW6RHQWfcknUNCq
49PHyyqnGFtcooujg6uyw8gt+v9nPtO068ocWslMEOdKB5J34YCJ5mSOUNFCg/XUsPYy/8a2ddRw
/jQTrsTgGPFkbiz4xiCgttX/PON53BU6Y0YX7Y75JKqiVRF+ZTVNZPoNUibDby//PxSSLHVu2qWS
fwm6Yjw9iCH/4Wj7DhmSAfxZRy6/HdXXfA4CD6AheGJ/iZEXq8jVVyphHD5xb2zu7lGi1QqfBfX2
y6hGn6lKAYmWSG+vR9ULFQXdTMfKEYNg1FjtIL/wZzEucrlhr3/68emPZpeneTUExWLeopToVEoa
XEGdSvibxlkoLpU/2a7DSuuu2c/u+c3bOusnRbmnbGE6nXks6DMNjYAfpDdxbp9HzHMOqhWifLoT
F+CzM79AcjkFWwLHRdsqnEEmVlkAjKn7PYh7LGqofFt7g2ewno7itMEJ24rR+9PfbN0MP8DXaXIP
0Uqzt8m73Jp7wUYlxYPxxEV1Ugax/J6+MOe8Dp5zIsaAkJynwUYvaN/B7RYroQrm37IDYJPVsFOp
hVx7dSBDNn9jhUmsO5uRwM1INOdakz6BNYxr7MuSEAh2qrdfhbK7hjHYzR65JoJx8GREC2FJc48w
MNXR6S1u6qdi7F3VEHjCumrASLPA3aD48sdpalfnRvx4bOFIvlo10l+NPzs6k3DCJ5kT955ybc5u
zVbaNd5JI2lSSMFpAlyfDPuj0qBTb+O9RX+3PvYNG6PCZN0BcnZle+P5SGIGf+rkTy+pRlVAxzMz
j//Pa9gKxhlged26epdWl6wLZzDTeWZtdKwGp7ZhlxOK+t8qD1gr1AXV6wLqzWOtDpDjgvpDqXRM
5zxT9VFZpMI6C/3PxZkgSXSnuNoOYiQykSnd7i2AOogqAhbXkRMo28MXYGYrqpdoGnwQIq7Ue6Vr
OG3Egy+aDkzgZAv94eSWgzZn7yFiePl+pQJcRjrmsTtU8Jt0S1D1qPTQjqqMSbiQS0+POx9o0AOf
WnCzT1WG+rO/orgAe7h3eysy5DqzKyPKQ+sK1+HC0GZ+vD1mJKIJ6pqb7xCCtTvrq5Ng/NocXWuT
87E+ZNUUVkg2ITkjYP/b2cezr5xmUDTBYepzNVd4mQ7i1pjX7eZvthKpeKxMIBBw88DNd/9wLicV
qGbnoW2S3ZI5HlKRBlsuqBGQMl23nVc43ASkh0gS8a3Ke1fpl2iMFlzNJgSYhG8MSAYZnb+e8erm
+E41loDXPYsRBdaTeYBOedE4S6UKInP3Xo+ygJWDaHcLq/0oXUTMlkIM7CJpMWRwgZ90C7XVXPYo
xsvbfqLQTADWuAC3hANqwIiSTKXb+qFHBMQHt9n2P+bvkMch3o+BMA2uYcJpdHYC/kbNmml7ypZH
PFZ+JS5ZUyF7jGEuklmtcRHrE6F4XjrCy7dB7wk/tJ7KY6ORW+okWt2x1rY9YPEykWe3zRTssAOL
ZLlHAZs0pIsNz2VOG74ZPnguBE+u+gOfZD1Si/DRlz8vk13UmBjymiuBNsNhggDFlpJcjlN+1ZkV
hMp2Hpr+Uk33tsqUKUnhAjTjoWR6euiYh8DGYzL070L5b/NN/Jappn/b8W+WjVJeJKO3exfrUj7a
5oe1iydISUmfo4RN/i1v35R7mPKz9n+JmqMQinKHXLlfOpVz2LU1DZQJn6UcK02+dJMNXUoRFVPt
B2264lrmochnzfCi/IhYnPLaSqiqF7ZIIqI9OniYCDm13iXik3U9+PcM2c2IEyqha7+Di9XMgIfh
1yOg1a+QkHjEt9jAXx+J3P+/IWUkX4qCaSRZyN4lppPoso/hLCnYUt83cJVrSf42Z2PSHaUFyiaS
/j8/nQ+Ug687qfEbIY2ymMEoAAdQtbO+kWSTDk+yeR03GR23FdeUdVsJdrddlV7//HxqaLUtdzhR
4ortVTZr+JhyqWCf7h45BvNkESgFMpnQ0DFTSoSYUYZ5d1VHg4aSoHldFazR0B+WNENnaLGzVsEq
QgrvR2hrRRrmNgeOoeqCVk2Q+2j5L7KL5WZAia8kRPaYw1emXfIhb2sR0xIl7tmqQOY6DWKpxX1G
3uyTdYX2U+17iVNqfbGqVV8MkSMOWC4woBvQTlAUzX0iacD985URgAk6V4yLBvL3EEYGMuUAUvGs
GrCP1wX5LjPMzRx2V8SlgGSOtvfXlZP4s1m5EPIL2Cqvojz04PJ+83MIY9mWPrwloz/Z8pwb72mY
ejDhAasTt7UgUHQ3OY0creKDbmQvfKgHB+w9sSqW5ThiBvHcj+7v4t/TUuKoQDeUkla6l1E/xB1i
trsHziBk889ZP9tGEyj7LPbiRYbPODe9wmsPRgfikE+J3WXGfn2OYr3LhFDBBuKvXq3808MRpx/A
832adr4JrhODxIJXXDlpIwNdoQFNZTSLwEDtIhCINWRSJmNGIx75ZPcFnlWJJHb0pVBQP55oZxZp
PS4gJ8of/+m2ow7iA221syh0I0lWWppCURsCy6iuEMHED+fkAMiH9Qx4ffSnJNrH7Ze+vyZGg4+z
z1biNwN84cfGq0zF5PcmhsT6mSNnx1iPKsVbPGonnoU9n6NJSVTIs5AZ8vziob7xaUPKx7AgAKwW
9WHjzI7EYvCjrI+WuDBpifIE0bHLzViZnyd8fW0BeKtRjsRbe73g8aF+fzh/oIvO1boWBVCr5wiW
D+xS84g3FekvIOsQ4jVYRsbD8L+PrMfwhKwaYAGTHSh2FeTbEwL0kNZu17Fdyo6Nwp7y6E+RnxJP
8vLgicnHCs8NPM1QLXJ90113XAohKWOkIqEgb9SItpVCLJpe8WTpy3txdB7LljekPItKF9gxJ+JQ
Ns3F/3ZEO0s7hRb229z6QrunWawooTzJjBIRN2KlxYosXvqDkUPotRhAmpjeELvO/zG1Ys8g2wjZ
ULKy35QFGYGVnkEEUHBIrIP7m7vyOcX+aSOcD/bVSMSwKyLYhRWhjIMdakOU+Qe0zAduQvmGMVZS
w8aBXlyPNT4cbNioqWvqkJQBMzYJoh9e3yzQbVFCQMV4cQ7C0IJ7cnDvzc2unhpmMz7GxRPeGEDf
yMSZ5yICAh04AGXE42W/zdPpGZx8/So1EatMvtuYYoY3gJ9qQGoF8fGBLVpcZJfMjMDhrIrzDuV1
X4VEYEZtDRBl8NgB5FwYMLBtBL5p1wapIXBzhvEXIi617sw40BC2JhwZYb/N8szaBVQ/vEhrjvDU
I1NrgONOUggKlqkw+GDaEK0RLCEq5Vmwci+TkJhCVzbn+60wRwOYIEEa1wTsFhby4nclC/ayJnX2
mhr1vP4su7Tyv7JsBxAvC6V3150Xutkc1Wl5KtkwmNzYT1nkLg9o+8Ta7DrYWCKZ4jUuU2p5mgje
4+7TSeFGQmJfIySOla9Q4Z3inLHZfeWSBIOAGrKzTAeVlhWRyyilLzgIoDz8E14RTliXFhQXN+s1
zYvU/+fPBZ7UF5PWa0fIRyMm//5CCPsMvDxdBI7LqXyHdC0U5ag4rNxzPdlMBJJQ/Z6sPMADRW2s
wyAytaFkX48nffwDqTxdR4vb/RoWNah6eGjTFNtz9yLoWMlTWiBzjBJcheMstTd441hKj3SJ0IPA
a1CYPEFJc40XFcw+NZzNQZvUdtvpX9txlLBc7AGPK0DiOffdycpTwGLH5C5H3NCanT1N2tmI8Rib
mXwnuVRHifHmgU0Djhosbf1amYShIsSz2bc1bVmlRGm6P/4OBMc0plPcjjOrLQQ8ja86xbv4QPPd
ncCv+Ry/Afw8iL3C9ER0NXouW+A6Lb1ikVc+5bfTvJP1h3T6Sr2mV5VFjNIYs6JhEpoaWlWWeuSS
0baT2KSh8McqDdWVQvfI136UjVAVdzQLjJiRRYqzKjJsxaOz4GwRHQO0lDUoMzMIXrHPSBqY0jGo
VqlCCGRji7CxZGUOL963r6SKin2Nvlyd2ofk+HqvqhMecGgt+4LmebgEyzahPGyZEYMD7XzC6tCp
YQu7M8DHyYYUUzeKagrGZYTB5jm78Zq/YgLBtQ3rg/N7RGE9nQclOmALkJThmwzGKWTlypw6zpe6
y91ef9dpn3PkM5KZH6uobigbqVnFtIwXlFU9ByuNKGAm7qY8zEpvopLx5Uujax7QLg2pM9/5WW80
G0xbr0/wFqRQnWBOODJv4vaorHgdbFdTCYknbg5S/vehABWjwjsuqwDi1pzQQTwYu+HmsZkclrSV
X9ex6KjoZXuwoIMIyaGagmu7w6SVGDwtsrCH5sEiA4fDiabrGy6+nAB/aXYK19MLxaTx1U8WedbG
W2ppY75ycNUUBinKPhEPxnz5O5FJ9TmFBiR8u9JMTMaUhNVf8uL26vlpdgrHqgv+xAc+hRY7Uebl
vM/BO5VZs4zW+5Gv5+DtBkImIWbPVbddKEwvo0QYabPXLPOcooxPrr18KrCzkeqWAmhGSKuYmYsy
HPrltp6KhWrGOlIi3cWRgpSx/nSKThElY9uGcjs0XxFfe+8r+z+9g5He4rSY+y2JsyquRqS6lTZp
GYBwDhePcnt/nbx51s2uWbkj1dDKUj8g64LK0Qn1TRIqt5d+Cv05nn8YNSU9c0PXKJ7hWy47heLu
T7jdx7nZ2MXZde1rdJcjuqR6NARNs3KTiSICgyuwYs6DL03D2zBGZa/oPjnJSWnRMcmi/VWQVefm
C+gt3BRrZQe/3LtcQJ0nst3tNqX4xadccJRh13/e1zR6RwLOKQsJqXFZVP4flB7UOs5lh4IUPB5k
GfzOjuLLq1dZsBVZCfXoFDcrQwTCTLgkCt4SahNQ0EONDvDYfmi3lztf1Oyu1BmPniVVkKynA5kx
mxn++o4xOVIkHFY6nEQl/egGYgNFub2svIXmfcCVPPMXtIygiXdw/b1KJw0xEf6kLD1+b9LnoQqh
nBkrqhTMNcHVYiIjPviZm+OTn0AiOwrSi0Xc52zLknSatooedg9qB6FC+ZgWFy0eF8oQJ+Ycr0ga
euLFvni83uipwKNDMUcVyXSg37aKYaNLTDVDlHL0hqjspHB0Y3c8ToKbCFlUwQzRpZZpV2nuy4ta
h/gWmvXhQln0TXBvt3Ro6ZVotPhvHwYjmmR/K01PKwMiiGg30c/h5JupE/Dx7D11j61sz+5d//3i
xbOokfjG7vfqSFtcQzMX2Zr5dhJbXucgDByy72J1eQLalcf63s3aqgQ9HccjrcAHzxmJMWIWekhn
P8lPAl0jzGCoD5ydK1Lxcx0jtcvN5bfGSzzw3oW7cIhUPFgytROSNtkF0rdb1cLBxBlk19mIdatX
BScafkzabbctSuG7eXXQOzykDOWbiVYZDBXZPKHZEzqWUCcAuFo6oJSK7HsGm0bVGIkCNL2uVTbe
VkdEduJUWeqWgXR0lbk9ldgQUixtqtJta+C5hs3C4NIpAqGncBL7QlzKCK5+ZgvM8bIzQHqNI06L
Tqvr9rQslZfoEumEvvRQGco0M+bPJAxbXWVrnHNGB4KgCv+ZTuhvWS05Wazh6kuASw7xs3pftg4f
M3djMj5Sk7lda5sbXqXVboMzZpOp8K32pd77fOpaGfNwL53K4XfLdYxicu4WMB+jwtLWrpiIaRLs
krMI4eOsgyrbJbfUHQ9WMpXzVu/aaBpjjHq35GDBaNtgilpDmPKxYgyksdy+WYFBe4iiabqNnWjs
xL59NjnWcop6PTf6oeUKMerYhOPj2g/Xg0KyrdFvBJ46Z9rYPWXDs9nmC3uyJEI5X2Eif4wjgUxK
69IiAuia+D1G/kLVmwP94MS7kfxiKiOUvNSIWjs9NE32NTrJLguVSCDzfPXAqphgR3v/pYIN+7We
LBsegMHj7qGoiqYOHhzqlS9ZykwHbEeEOZqg4cK1fTg9qfCStNzcJVwASp9xEWh6fhaBT1S4qx/g
FFc/H+dUlNvM0k7RIG4rwpnnNmglI53v9CZjLCOkpN8w9PwD6Hr57UI9qjMlqoytJ5J0RBtgLlC7
KoMPUMHeNFbmrGeDSzwoYje0BisnQUhn1eKgjRImS7SKyjsqQBjjxJYd9eh7QGMgxxFu7NvBfBef
lWsLaj7B9afu9OCc6wJ1tBrhqMs3D60fk2qliS6yJrtRJxz7NBu15UiYFKuefvdybzfY6LZFB792
09ZjUPpQ1PbYXlM287hM0CTmatF+JfKZTUr3F587kQdQfDnOiBsaoF3La9vapzHaQV4UEGTvDnW8
rfV/flGzab+9eOBPdhKTQGh9xyF0ZvayHM3R4vR9RZKVOdRXtqzT5SwR33lvSVbRBU8gNjap5ML8
ZfoUO8JyIvXXkrbxJWGOYT24IdtmLVEZ26SlJKYDoCUrNsf5eq7jD14dRIX3dFoqtu23LsthK9JC
dSY6pZM2HJUWkgPvmf2QPYlL9xwnqkQNV8jBqsiacpaqAi0BXgNj82LChx6qhSNQpG4EMDU6ClhR
4Hui/XfhxxBODTucEk1dytuky1ZVfFL6rvsSGQTQBiR9JUZzrbsIHGHEe6nmVEVWmaA1tMKyXZWr
UUt1W7s/Nve8a7ffKuK+vaIIAjz1Ft/0Mt8H0Ey3RvrzLN2l7NO0fDuwyduDGIMRCsOGMTTWqyof
1HveHXtfDfhmwcSao2FeNKH3XfFVqeIQSUIFydMmaBwKlGkAxS/R/IN1CDG5Z1LRH3axvUEctCD4
BiYkYAYkxcEq+mGrr8hkypMHHjVhIJ3I902P8X9yWTugrUvizdDTL3oOYihmhlObt4VCbeX5V286
p1iy26GVSk8VdH3fT1syUtt8rNyw7UTUUi8YOZO1NKIyu6nnCjUgCJpHURbfX8cnWsxL412Holni
7Swu4bhX3yQw5AIbm6XzYozB0sssqRUtWWwe25HZBblwnUSooRWaBEADQUG7QfKfI/d++naUkEWV
FwQwn6glRaGLaRQj0LDLZUsSxY701U/+Z9QWKuKE3h0H9Hel0ztr7oeu4B3//qXhRW9LOieVMsHa
AnzyUGaZGWMDessg9NGDD2fKPUax5MvrAiqS4IKx98BbMzifBLSrQwgLNMjMDowniSbwMeCrfq1G
IfJdnzY3vxB7Nv98IrTKVUfe3zAckkRectGU9RmqI8qI2H1WQ9oa/Ne2U2X255c3RTT6fLTjbiun
2gw5r5C23s47IawxVHVaLJsfjb+kQUTCoOUc9ZtDvzPoiQsM5tfMo7dyuKxQsesYdZ8AKzBlXqYf
14rC/pRm/mwmChAfxktk+HGTEPtDJvEniymS0sDWb1N8NwxeqXok5rdOm3xL5tZLmj5e6k8zKOkX
HMmGCste56zqyQaFZCSLxyWnapj4NCyfXfCH8fO1cFqgJB227ouFpMBE0iUfEY10b6KEN0jbjjrL
ECk8xgji1GF5UUGnAimmJBOlotI9HU4SaYQXVNXU5FDBEZEXv1bKOQ57exj8K8z9J/hTlrYvh0Sy
utE+xEsa5nLuysdpzNQJx9rDE12MlRpRAxZK9DZuopJmaqTo0ZvQARvvIXiQ7zTS+ywL4B+hzJQ4
Xw4vaH9idxZwxU9T4gAHPfr0eNFwjFsEYnH+5Qph0TIlRvGf59nLp777VVqGCGLgMfQjCt6D+DVU
3IYQVI503olUKQt3c4Xv6v+9igggqLB1Gyf8EyIBPY4QHDJig978yVJPprdKM0GZ6k+LjQYqJtGg
iVNBAXWXWdGsXT0swXcsiCRduiR35unztMfem/9h5coJBWw0FRB/XSBZF3msqLSz55OMcQTUbt1n
PT8mKvmAhujYDtoi5CbLRWG7FvQRDug8IYGHa2i791KfFk+xP9fpJR/OyHXGduPc5gDAMjN7eN+q
A45BlHo0xc9SiAUcg3URmmzi1wHLgWDKfkA1LNvOtVweIqeEsC79QFwFt7XGCDKL9Iu6TryvZUTc
8IHTY3iIast+GY2wlnNAegLT+IkFLvRxMtLtt3/F9nTntyQmDT13c5rIofDmG3y+CIhq5LnioMEz
FTxsrHTlqWHwLtVV2HeYuOe9vSv0FqdqqnS4dKh1/VH1se2ouHWJXOSM28V6DRrTDsuaQBbjj5Ia
R8m0WlnjK2cUFsRDwb9fcBDhxAJk6O7LhoWJK0ges74p81EkMegHLWEvqkUoRhvIjCy4iV1nUjPK
FZvLiigjMWDaMV5zA97hGdWLR7fRTqILtKGnJzQKl60KcSVGOCWEXupxKVRGmTp546OTZYZ7ttG1
Ta97PD25nr7N9JfpweIk3Ld6LrPIfY1I1nTM3BJsHITscsvl1puxlFOErIrhaZkN33HImwDlu3Gp
sTKSYfkgYG7X02O3t8WdmF5dArrUAWxaraYbbwz1f2vcUqjJQbLb+UB6LfIODhqpql3NY+Wn1JLK
9QCIyv4WX6pBKXpQnLJeUrUvHtrkElJYf69MxJtGJ2SSjC6w2XrZLJjWtDJ3cx/3crHUVSWYsg8n
dWjt1fsy2gOrDj2AR/glNG1tNc84ixgQIk2S5qw2qn6nBQNct9J6OoBKMkYIXRjk6oDUzM+mh3RC
lW0Rhd/B+umilFqWrpKFMLS7dKY4AhDPCK8an3vpkT025M9qUOJzzHg3hp7u36ZYzsXks6LsfF1Q
ECY5CXqZcKnM52eYPo9WdAB5X6GZbYqs2vQdX2s5ek/uopBpmN5yjaQUwyfBeEZkYZeoFdUao9am
SalhUA69qYV+LlC4Q5YCOrvW6CDnTDogv2sQmUj/mq4WIYVJ29vKH9p0O/G/qjQUSOt98eYEPlxT
ci+I1yLHYIqPE9YvxhfmHX3MAmQ6SiuCayoSoxVlP013Szei8SAkLbj+nyNOeNVx5JtR0qwLpeqH
fTS/TxCeNQbEQutBT4ilRe7oHlmfmGKKU71H3c68WuOlxp8XK0blyhB7fmL2BhSBY7Sp+A1Jb4fy
1v6BaDQBNsEW57wZ+0nuAxvNM3MexU791jHaNOEjikqLlMc6tVkn/864C9Th6zb27eZd1T7LTMVL
Mup5hBW3RE7QaOc66cmwnifRLzhwdWG+6T2+tq8vkcQlSEaFsTWNDBw+VrySSmQhNmVnEB4naiwQ
bzz3qIFZfEasxA5IvkQQyx7GEHyqOhR5RVuIZ8hG32u1Gal4yWGoBbiDCdAYPHfmFbRkZIbovkeP
+ANo+sY1/oWsq60e/bCumo0hYsjItS7Mo1jdAaSt662lwQW/Ic7mJrvLuO6Ewwd6QzYmMfFkgAa8
WLAgRY4BOyYC2wMjYM4XR7tYZ3w5kvJE8fnZhIQTEwwxG2ViT2obWOx66Si7spC4YQrHBmDB9/7r
S3vziut1pGX1HUZUThzXtHctG+mFYWAVjL7+SXlw2hiFmRMqEhvazV0Y07YZ6P8ocRm2hmBw/p7Z
r2xAa38dg5UhwcOTP2PlvCIdFB49vRSc+HvQe4GMqrM1ItvE3SMJnrAIvZQ2bA90GXdp1MnjQA5x
GKXvLPOUTBIIzbEBEClmzlDvIXD6UPzh5ZlYmoR8TLYBIG2297iYX03uTyv3ideyHnrMcBLa6ANC
a4IH+sYaHH7JBx70RH5f4zsQ2N7mmz4FLN70no5CDK9L3cc0WXAdp6TrrhxxMhIB6DlvBVyA2Ol6
HdLya6IUSBTcTSSecx7ZP4JKPD3en2h3dj0mBtTH9LdT6NR9fVu6Va4R0Gh7X8Fc08WD691A7B8D
M0q3VfpeFN6IgBZ/3MXdojJwM+OqAoi3/b10z3fFjeIrjSsCMsbpFgDt5eDTFn0+0b1gLuY+7kYg
SVZh4Iqn7oxTkaTzNW+YItR/bOD+JfKhGK+N9cgvLpM2BkZRkpeqjDHEIG2pstY7RFnS+Zm5Oz+z
wBDwQ8Mejgs6UpY4k9Z1hfXtIIeVcQx0aVvNrbdGMvOqIXCRYz35lrGsEAOY1GLBEfHarogqFfw5
MnVwgzVMUqhIiDz8PTP+vVls0uJGrg2wHy3q1ZsnUvouGLlLWA2i3v/G23vT1tvTcb5p+cMPbERz
I/ItzvWi+PinJiKZklI64B0/1yCaSK+gEgEbWdJOwtXZDkVAoXlLuqCyGg4KJ+EcBMscWrcTTWVy
bZ+qEMLCo+yJ3vMRUI+4xwf66s+fIIyPFAnsjrpC6ea5uYy8pFY9TN0dQkjpdtB+SRzLPf0tN9Oy
b5aSqDTQBdex9Hd3y9z1Ysdb6HmsQhbfjQWfi2hZmgJhBx8X9MElnLJKaqjAFE3Blfio2WUo0nAr
jR+SREy/7a+Y3FO4Nu3v6wg+7yg+GXxFt3uRCBd7irsvViq4+nc3+3AsjMfRuYjNiJQ03QN+Atbo
RUYF0RMhAJ4XHyNwfj4DeT7lpKfgEIGF/qyTaGnHZf6JFbNsOeA3GmQp88Xc8bK90cwfNNhdkfrJ
O+oHCkvrO3ais+0PLwPLRfGUf0it0vLkZiy/USz6ncLM+Mk5Ble8uJwZHa/1ILMAFVJcDje47wr1
O8WprhYXhuASTNdwOrX9Z97yEVq/g6nh7ruFQy8vEtoTRw3HMdWLDyRYKJehTbtZHK6QHyOQ4w8w
cSVHyxo7HurbLB6GmRwcx3VI6q8Vcmz5TDIgVePmUAYyt7maNlK4iu5TTQ7fLm5totwSQfyjqOtm
BBfr6F5hQjGvvJwVLn7xQoRdNDFjNRvpDOhr6Bww5ppdTYhQQfZ3bCvDNc+HMcbXVHDkVRMsBPMu
+1+jxYmHjyBNSzZGTVHfUQ5fFCNuZ/qbvtoDqsrpCzlpkV3jZvHpvrWNxSJMQCHVyBLNqKiF4Xqu
ApS/9n/2dmb5ROq/CABmJfsyYMkMBK0hb8N70X4F6ioKq9639KEJNkwnsX2FIVG/uqzGfx2Pj/vk
FCrT8xhYeJCXDIDkwJgjfEnwKXXDefc16R+m/KmSiMzlneRz8oKcu220LF1tJ127l3R+oqzYHuUz
99jRFPM4XmyDu/Oq5VzjPoYB53LyjNgJOj5zSRYoUTLV90XlZj7UCa9hnjNjsAWABeUiuvUX2YVy
BWc+e1Xx1T7TJO5UKM7yPUl0cs5EgmXfrDtcbU82DP5qca2IelZVbEdgNW99NhAm55mw6lqz7vn9
7iDix/6vvVkgmWrDkHiHEYLQ0HweSfg1dzJqYMk/pZh5ft2752ZkxBjGweXBjfzB33InXZ0bW8rQ
H5sOYAlJ2K7fEKd4xm7JrdUTRVthbd2D/EJaOntAYNyWktF7sdfu3VDjwiQS/iIInTp1iVBbn00h
MZ7EZadF24NB+1Vj2/1MKw34CCOb0lpE14bAqAMwtQw+wRyh+e/3iQLdrYmXi969bJcx3VOQVybF
OvyCVbszArAbkc/BxLN43uZFX7aOTfjFnR5w7ks/2lMfrn1nnsNTFbe4Lcgnhz5EB03VreqaCium
uJkP6BwzVrv5mys8eYy0/rhx2urJx1EsgCSICc1pxnJ803SmUy3qKA2J9yJzL8kRu7CvjdC0As2S
jwhyXBla9ikcuvMCmAVhXQlTO2wqR4l/+rrLaFxAPAq8gtBTcU3RGy4XEN4R+SuJ1NiMeeKm58ZC
8EVUdG3PJ/XeRzD6oDUlCxNSL5nz2bXRfdtwipawHz+qIyHaKgpo9WbFpSMLm1Ywi/8fJLjF3bPk
J++uQI6g5/38yL1ICVthXpDVAHb7UjoR281exC0ejY3rcsJQmXxbPGzOfcLimDyjmvoEHR40prnS
4Xln0rwJC0EtMfN3YrCOYZxNKsMVvgUbUVDPor5borbQ3wfRnVbMd/EnCo8Hq0r0/64uLJfzB9u7
csXpZ8SzRaXlpBOVGtUE88pMA1lPFJuAdxDk9YiE6dR6QPwgj9qftnhyTC5BJwktZFFQssG4RuPh
DcZatfIdwLxEFvjod2uOMx7WeYpJVCrylYwbKXxD0WIqSs2Si8l+5UJuzoPB8jFWaVqT7BVm4hNj
eanGiHiyPPzKdnxZrFfE4uauMU1UbTdt/wMvIEAnkpUYsGlU4NNpJz7Ot8IjA/NsYx5ovkSrpjzC
jFzSt3ekjjI4eZTrB6P7ExvsoBS/ZWHGI1UHSM163h0PlzO+W9C5WYopXjn+flEW/ALmVZ38nGwD
ghEehJnyzhJbCmo/vX9VSiM0wboAM1Q0PuDRtUaw2T6qZgQhPAmC0ImkGsyYdEAjeCAqXR2RrrVy
hZne64sYLBBiZIk9bR9LIw7UVk+GWDWL4sKX1nQ4YbavoqtngMoXyGuDZRWiVCGnzioQz1Esm8e2
sFT9qR4SbDfKCGlZA/UnbOOqO0RHjH0Ishj4sUDvUBSndHhFVLcai227hC12AD1kobYIvJj/jXF/
m2SkOKXnprEQ0d9FWnHiBkMuj56pndplj56cAcxfXJXiRAMBKBpuRB/GEMRzZloZNdRB9SYELr9r
WdSPlOHouwm0B7os91QwW4dUXe1KF4KezfuNQGzZG1g3MEYp2xzWF/uVUZQJcXQptLYW44+a8CaP
l2vHiYo0oasODV2OTRcCfhtsAw+GOKfnQgvDOfgHs4tLjMjE+bWvfC/JdgYAcAvs2h1AjCwCUTox
mkzvXhNXlYSn49/DwntEcIG8/udD2p5IXsDLNO9nqGnaKq87267tJhEVvr9v6R7ep+7ZAIETCDcj
w0khXGWHLeol9G1J54XuZ4TRi5Tyzh8D46d7Ar7Doy6zPodIsQe1OTHm3PXEoK6/Co94V3mnqH6X
jp6g5x65rhhpGmA3VYmv2q5X/No+3OA/wF8QN9l4LTeU2OxlcVeDK5vMRI2RoPABvlsAHyUL6uti
PZJ9l6qEkWxgH9uPX7FW2LbYvrUocjTsKT/I8W6qEzUpzRbLL8qpZN/zBTeMQhso63/YMZpvsbu0
jR8iDJBBBICtdioEZDGFADjHD/pE6wwp4a2z+2JcriysrB4e1Qc/HGBvkl/DE1L2NIVfYqENcxAX
KerY5mSZoXwMzcDdkmYrwJMjL8PNdRbMiUJSJtiLv9vJIDffDw7Z4uZjwWQyMr0zq6ZKJyfz2sGM
EmWIpKfFp1Q8g+QrvplwnH2kuhoUIrDiLkiOQCvPF7DuwHpULGpwpU7CWDfbs5O7yhfH/Cv9mTCw
/A6zKMlKCBKuFmyZXkWRzT8pwNARPRIA30xypNcyf9CVmQGjEBrp91x86W2WJXNIGNcAhZ8MkRSb
46G9wrRnNzoELowrsQmYb/IDJSSGlcK/au2V1MG2Z/oWrGmJhaSv2kcqaxe/JXyZagk04CNsf0Py
plT+ldXmfI6AEnDTUaR1cYEpL8U6ZPVyuYtKtjLXz6QlOF+6HbUhlkEfJMrY5IfXX4P21R4HiNXM
1NeaMynXYheWHJCW+ZA0VI+5B2jDkHqR01LGwiQ3BPyDKJ6t9kf4j2ARZP7wfTIlCP2Fbhea5NIj
HF2siYaaZNqikTjFIi8iMkk6BXrSl9rFmHF+tvpuMvs9F2jw1qMnF8c4FwqGVCU+6T92IgF+ie8A
bsfpBuN6LhfenwvZv63nOqpFNmFAfQvTcKc8efkTVraQZjX8pAJoMBR60mR34z4O8ybB5CG+Q441
faaBWbtUChCHX0IlJF95Rku3k53RfSNwmLvcR4AKiA5yTHDEPzLQNIk0N9tGHUir7uoMPFREecOS
E2XmfFhSaxzMFv0qZkkyCYNsGoSRdHjJXlHDml+1QAScgqMj06jihcbGPi/se0RaGlAqXGd5WASH
u5TjzRzO9euPHwhxJxr4XUhA9UOoFw5GLegvcjbro0Zz3V5S7nj2/mgrKUWavpmKawo8UnS7Zm/t
Tnse8Rl7Z2g3rFjH5rCTQyPgdwZWusPVdKpq8HJCYtFTM3cSUDzVdwij7/A3YdFwSva0J4++zCtU
erqB06NAlpcrupOvH2tJqT9Dn6qNfks9xa2MFL4fLRgeWVVJXAupwCDQuo0dQlywUee41JjNwAIj
LM3AWfL8LiwdIq/FRRcJSLtpAyeU3Pltb3QzAwrK4DbS+SBOwBsg8nmmb98iMnppwGlGkG5nzkUs
U24WpYOHLW63XWU3VoQCVnyIFyPdaFicQiIE8urBA74jSQczgV5KDlYXd+jellVjN8Xr9TO0goQ4
Z2d6rzQG6LBjJn4dvHdVyzc7+EVEfAnZKyr8EguQuHREHp+ZOFnuPnJjgdCg3Jl4Gw1Wpc/PBTSG
Yb8wnpJNKoXLACcIEJPuPRGLwMF5HdCDE0VGw7Rx4Cg9cUX0SHtos4ElROafNPq64sBvkXm6JBce
7FJN5i+dxcy84i1utHHi5URdfx1GWULmMVt8FMmOhyDftLUm0JZUfpUKVkQdee4KCDRhByMA+nwS
c4yxOHofKPA1H415IQBBr+B+t2rMCwhRCWwPhYq8qFFP7YUsdwuS1GHCxGuusfvgMiMFxIhYNn4V
PvL6wU1AwSrstWDDKLG4130eatISId7xcU24M28JYqbuGgEhL8us5USfD8XJDzdhHagxiMZgoyau
YUUfZTrNASkidhsxcNIYKnXj7ZeBf+MksANsrl+LW65hyZoqW9EoYkM/16m29u6dLiNwXXaI3/Ew
8Lm8HixGReq9QuJKLTbc76ykMZzIOwyqmZiseUPFlfUwp8c3CAu67fwqG2Fxl2HK32uws84c3yE3
Jf2slthmsbbm28wS27YPxG/zi8Yya5rSmgBD5i+bH3ZjhT6keFJ8LJ57Ayu6oKH7Uh0HkOffrZQy
T6wNPjDy/f3YIwpKWUbkq/lfqiNjFVRGIbMn+26btJ1ZTnvugkLCRJUI9DY6G9IeOMxDvx+Rp0Od
W8Ji6475zo95eh3Z72zIQoSgDas+ikD5EpHe8UAVNMEoWuiApQD+Lm67tZHUzMrBOmHCnbI8CMlO
9av4u0z6xMji1YeUKSzvXzveW6QscMzJ/8Bo7/sD54PKYD4QW7nkDuvFgTQyjx5pyD/KIim7u7nZ
A+jDre0M2G7ONuuzBYfW0CyhBnO9Cl4PJ31AcY0rOREeCr935aUcNJDFF5Nr47k92xfH1GUaZS92
451GLLcv12uZ5U1HsimaqVZKkLHE4Lzxt6Apytd94DlGLbAQRj80f0NR5dH+QC4Kt7yN63GBe5dK
v7l3AWJd+lfSBAkDlrND/wDTSH+eif/SG2HW79WkDWidD8O9ALfMiG0mjXdxVX+7Oobi8CInfYeD
DF81D6SaOuPUgWA7FfysEmhz1c9b1nHSmDuBJXeKdjH57/xB8e2GHuyYmg6XZ7T5pvlpqo+cC+qb
QNUzrM8HciW2MKcoKvvWQ7/b6Ksqcr9AT59CN7au5QuHpBmNmp0vHPtgOMUicyMuN3badHXJIOvY
dIjri229xLOIqIn8qKv5maCTke8A822EgL3KoKEVvQaauyOyxGQvxDaFMV9YrA95G+7kXTzfPF6S
4ZiiYax5XXPJ+y+5TC8tpT3wvQGJdyrxPFG37BsnClb+CnnEmhhJu7FXGhxjJ3TAdxCVrdOgy7xj
1Q+futcyqXbp2SD5rIm8KBz66e+6y+ZnTLNmcZ0Pdcx8z4WPZXSUVEdhfkDpP2HSORPa8dASvyrw
BSpdy47mMyGe3VgEQWaskzAzQfiEshU7DNlMJUIHMKm4TkMvzL6tOlBJ+9t8vHOp1TUvbZB96mTw
kqfCnoeA1MglcTVk0Xh4Q759KxG421Ggsu0Q+XjN4JjwY5JWDVZ4yWcyB19C9tZhLUSGSK2JtiOI
Xxs+/OliEjkIi4sXYxYcAx83nZq1EhABSR5DjE8S/x2l83VWHFs9q82hUj3U5waQKTz3aHob7AJy
alAFC7RawqchxkfIivY/Uzk6h1EKH55nQx246qLtKSX9b6/j1dNTc5km3GGoA77xrPFN/an/uQmJ
lJYvSEPuIqBuzFO2ss6jN4eI0yKgRRIb/lCSL+EtnUJZtqiBaWdyUG7eNQTGIG+AyP8h06ujYIky
HdKOWGrayHFpmBwOgUcF/HbGjd1Qzgh4AZF2sggQz6XGVhTVjWa+IsVfN1fYM8ftxZz53Ysg6eKW
crbHx54bcPq7CNjXTaOVPTP2/oHk7Tw60SDZ//6Xafvlxa5xif+uHWK8bahXmg8shqKgrUWH4HvK
luUsTqEewe+oNTWiRVPtqhLHCk9ZYuz8nnIKBNR9yyhwnJXkU1Sc3XT2jDvk60iZ2ZEymPAnxH48
w/lXRmmWM5gDCIPGAF94WA4UY4qXmv4Bkul+LiBojH37+l1EVKFxSUNfVOVTbzEu6Zsqj4jqbVeW
qyg8FjLoSxKJz6ggkCyN/Ec1QaXzcndYXfDIkl+bpWSxaoxGwqE1tr2imJ7dlAcsSqz9EyW3rVyq
/KzXguS4uUpmKqCnCoy2POGJKVS95aeki3uVwtiJx9WPTmn4cVLRlgyd2sUrWm0HGAvom9RCShhp
y5fEanoFwrcDb+foWn7a0onxmiGVuLMcZZcGxrbj0OhNuHdMME/ZSkxqS2LbG1JE/gCYWzXCQ/NQ
iHKUQplE1re33CtoHs5Ascvcr8g3d8TO+bHUV/YT3NPE8avDDCJihk+4erwYG0YSqq5AJ4/BRTaj
2ytcxy9i/jdG9Mj6MhIS+CyG9SkupEIhNShiwkyjeSHQi8ifXfzwxWlQz8698hWpfh66Hp4zkSmG
T41bOqGHax1pmtS9KLMV2kQKc2QOqe5dSy+GJ0zxffC4ALJQo3r+X7eWdIOdIpZ4VCncheX2bf/a
vfQLib6Q40r7QERKa/dllPN4jeQy8Vt1XVwbTbiXLqDB7KcLf/F8k1yK806ItesmujIhGbYTQHFz
8H4aNvYsDXCPi9keh304CHxLASz8BS07LBimGMD1tW2g6gjzZ6yThrSE+YseYKuio13qJqyA+Xhc
LUm5zSH3wqY8uKjHSv81QymRywA6pBgmjxQO1V0T9eBL+9kHVvCVFzMSIvS+NCcIq3zDl6htmJaY
lqcrxi1sr9ScvOjssk/NhELJ2tRxZqsO+8ZQ+D00zE58PkwCc6tRi7WtcLm9qLseltJojAUAoEB9
G6FYx4fDZKKmBtzpWSozRu/QgnqsfxLfMHn84qT/Iup4xqMYchiJ4x/N3nIyE4CX/+AJpqal5Kn8
n/V20NnlNs4xoz8fiuaAqLEqkmULJvXzBr7QPz0gcrux4plVi/fCIDhKSX/oBUFP8ofBAleLa4rd
1Wt/VuIWJBB8UvVG7jALhOyUXXdQUvZfjGKW/mun3NBkb588ihXrKS4FXGi4OkSvJ3ETCvKWl+Tq
lqgN6HYYkeIcL6+ItYngmiPbpkCrAuiis2VepnYI+iR789RYuSkVjWiN+a+gXho5KYAp6m66NIXN
NYA16gF+c5+F69i/vKZq4fcZ8lzedoxlKFafYrjSpq+E2ynANd7NQGnLNTrDV/TkUUeQ67IovEuH
LlpPT0Me9Afy87yB1GzQ1zBjLdeAlvM0sp5WFK6FvXYonIt+sWfOlJUncIuWOJOt26DoF3Agh0Np
2K+KkUXFRxR1lvdP3hW0t/9MeKq4Rjc1Ey5YG12UwWTW63hxg51h0V44ROrSz4c57YzQdABMqYTk
ozNvDpXX/7BA/HxLaGfekp+eIz0CdpvcGumi9IqVAHOv8Rflaqdot+wBBdEYdKXpd81sSNM31InX
fVq37LRyUJ5bllQlyrgNpJQru/HEzn/Ku2QTxIG7AgRsX2prSgoi1Hn6A2DyQg0d3ad9y+Mp9jhs
74KugdMf24yKPDztX/wgBcMK7GhhgXgKhTM80lowc7batNDtlXpBep1JOfy0DiTNp3wCMZDdvicu
zygvL0zs1OFgeg2XvkDFLnzIOwtm9GI+457el2R0IQxY4Rvk9PMLOsVnxwkpPtNEVFfxFc44kM8x
tOa9Pq6htepnnbwmmCsazLwas2eZTBe7ZEubLhqLTAF45GY29hPjAIak/ACTK1Qk6KHhDONGufu+
W1xBU1NXlJHT9RG+OxJC7ExBGAgQ3EHErT4FgBkY6FoFTEPFkdZ68a0ho0Iq4R4N979JDrKMI/VQ
09xS37v7Q6unEn/4hCrrmUXbLe+gYM4+WQNIWtItd5iqH0K0oCQCn5rIvaJTxIUkSH2lC8FaWu36
5v+S0d3E6swzoqZ5s/PoYTVfI1UR2+fWzQWo8DLUBjHpxenbx20tOOp+haRq3HDhy7obzlJs0bg1
3DteLHfQYJGuVGQIXWPCEnNWnnVQoL6bm40+AxUsbh2TQZa4AZq7YJ3mwvjSo3rnTnIgE/NfaeIe
NN/OfoKlB+3AByqkAXWNdzVJIXeWObHQwERfgqEvrQssVrDDL6sw2q57jNJhaWuPOtBZi8H2sl+I
NA0TRg+ERPJRfdtsj8Klqu0RrPFTmv+BSXQpDBYSTHcEWTF9yeiYRq2BxAvd4zurOpq0EXtR6CMg
PAhb3H1pXuEMRaXk4sud+qaCe4UTPzoV8cFx7ndqFC7guNrnPs7xmFG5UhgFNqT3Iu+QgXncYr6c
2EA1Of1sEQNsyc+yE2HUSaGbHqa5QCXyBX/xsquMophdQp2GYHrt6KI72zuHWcI1jKmTA0P7roB9
69wZqrC4uG8w09SkMgLr15HMlhhmaNNsnhblIxLFGsECRe374CIwxGgSJqNbpR8Q+fxWVZ/tta6w
DQSvpknhN1YVp2y/M2Iq7az4xWd+4Cwi+FvDXG223/Huobk1t5od1W9h773HPbUf/RIDDIOYB8VU
wAVt2LxM4sexkfZ1LgwR2aREo5g9G42kB9eFhjMmVFa1iybpaScPyt7L9dcHZqQuwNOtMVhT/gz3
8fTOXS04B26Uwg4HcwoQowxO2VjV5ywDTANGmpDNHYNI9vCG9tqnucojRjNcL23AHwGzTu2uUCmz
mu/cu5CetuA1qtvFCVCDbJ+Pf8qLy47m05PtWSzz9RWYCHySE7xWXzzZyiFLr39F1DCfMpkwAZnW
86OQCRu+fAkaTWrVYXjxULQc8ZLaoJQpft4fJ7WaX960vJdSA7JzSEwaamLWKahtHJ+T2oeOcH4G
ZN33GdhC+3q+f6CPi2qLoZ41VZ7buJDVQDd3tBldnGPcg2bQvLAz8Eg9FYC9yhGP+BchGp8J9eo5
xCza9GeMMbGGZJ5WrPoAyvYmQ1V2qUuqgK2l72uk0yCV3K9svcXe3uS5geXgqn7PC7k/ETA+y/E5
D3bhbP+zas0XnZyA/FQwBmJxmjBVYasuhi91tHvjlqBZ40AyM2cFGNRhucchA4BTckGuiBt6wNCQ
tNdDrQHMELy1sdXwC2srAKCACkg53wSL9KoRDiQY5owZpIi8Mfy7s0Az9ZXmFrWwOr+srAGOAg2f
Zwpk3+f1OLNrBQ00gb2IF4QDvP2HmyDZPvf+/o+3BOD1d2j6h4N4yMMQEfDaIF+vIVoYhJ/L3Uy1
xoGPevKc1D94vPmKB8XBygqpf/kxo/3sXEJ7Mo2/N7XAHPEoAJgKBTmuoww9TfRLFyYbjaO1LneW
51Src7REWN654NL9HWCcUMFhahf3EtBd7gDX922vh9fmqsi7kH1aARo19eIVKc1+2FbELXMgliPq
/X5xZxuLCdzO9VUJj2WGT1MRy5NZavCqE/Un4YbJi9g3mGTolM6PUc+5u3hcypT1Dc8+11uK+AGc
eWr8pbdj3XsYJVmaJnMm2Jsm531aEo/Cf2fKu/aLtpgfOwrBGjgsoi67Nibyk6DSUcmMDhYlTpQj
QhjOUEJG+6VwdXw60vfZ4SqwGv2uo7I+M9zTUkfxzdeZYUdT0ZNL8XzeZCe/xVljQ1ivgZmTLMdC
g2Z/ECIcxTPYh8ycTvpYCrjpyKNp1Kx71H0YjcYOzvKA70uF2Av8qn8UmPkhfx2Oct3B8Ggh169J
qrA0EPI8JKiqxmUktf64NaXBDFl8ARkB4ClNtF/+Tl0MTNbZDEE3axhfHJI2U2CWg6YXhPfXhuVq
KYEYfBXeUSVOHHVfH7FRiVKIbnbM0puc3LVC1rZ/PPWl6S6vaPT7O2DQuT9nnvn4ygF1HNXx1G01
k1D4xAMQgWRKSewX/bZX2CnAOrSsa8uYr/u/77SXbsk2h8M3WGwA+Kvo4tCFFQFgT+pU2eS/9F0H
B9UawMN9JJVz74NPrFQ0f34KjRwpDA85L5FUeCbNfFVDjir5v6+nQqfVuGP5nB1F9wEOOHuVAVdz
/5pW+AoDU2tx261/iZuopVuvfugByf/aKhgnYTFY8+kj/oQ3yPol24TbNYB/ivtT/zhFqhe//aDw
LP56aEEnx2FQ86OKGvTblGv/Ubt7AtrQVuHjVOhpcykwNR8NPOWzE1amtiCXXmGb1nXBJtQsWEwH
wD6E3NdlvOODHMiIUqocfJSiyf1n18TIEpwkyX7zq8uzUdKef+fEUv8wj++Xgnn9VuKGNAF4TY+q
J5dbL2fT6FvRmzfD7bdUtLu3GLSnQxmySwR/FB0m6XZa1v5i08756ALqTz+bSzMX00hZuY2s7gn0
9ohsLFxADpjNMuoyxKRG/BWtICDluEn14nhoE9k4bF18MC4SOD0ygcGBzmsLu2VrYPnGWUP2JdZ7
CiVfoHMlGDOUGUnjFt1hjT3YShhVj+2zLQ+j0c+wn4kmu1jJwTIiCRF/Y0erNJszwng5L2grPioe
rRJPrFxtk3wDJSPg7JGxxjd+wq8snI+Q/NSRSmY2Wu/HOTuQQEJyzVknnhwZngD0Hb+awVGg81ze
WQA3I2Mu03wNpGGAlW/dGJikNxAXaVCjOkvHzRFrISjHOzR/Io7mnR13DDWW1jRCYO895vA2a3q9
1CWN69fQWppBtYV8mgvPEqWeQLnwRYVVuiMB2UnAI77GkCiAGlomooAFYWNB7l/FX7/x4d5YZxU2
bqQIQc9Pi9ahK2UKhgMcJbcvsxH91xlg4FfbA2ROtKJu/B3lIuKpMIDPW5qxg6EtwEC7BnHmpOIw
4dKAe8rZ5xWyTSViSvDTmTzFt7BmROT8scBbmLrKvJQlLBs1VFT++8EjeobOF9pK1CFzpvEW8Dxa
Znhh18WK7pTCt+tOqMllEYftCqnl+7q4Um8eDGspNb2pPcPHe62ZrCn070VkvJLYljuKbVAoWFfC
YDc1uaSgOkVWRIGIciczM8byOmHOu09fMPEEg8sF3mswmS0kFnH1qulC5X/WWXbfjogCNQAAsipu
5357WZO33J8sZMHRxBSPKcY6Cxz9a9Q5UZkEDNxjsmWOBtrG1QY5UMIA5al3hFoQPVvRRn89XF+s
p1WGC//uz8TUt4BWr5QUbKT9XkyQxWAVXGR7mGygHStpDa5SXslbf7s92kjyHuFqvjwKtgBQAIQC
cMmIt4KDzAzGsEwp6ZhalUMsUBA/fWhPGE8940XvSIHE3evbiI7pbGHK6IEk/UtoMFrk1qRs4wYn
asRznsr0lu+93VBvNZfgGcxq1eSp9HnL3pmc4CVm02m+fhDr9VZ2R3EN+FiLxQZjaWAvYKJ5m5G/
HELS29YMDMr9Mw/UWPvFzPc3TnnUD9az9Ggoa8FUNb5OHeWGLM7lFDJqHYhuLTcSOCE2DnJBibri
3LDuoU+VkaRdwBoY9XIoDc+fxCjtvQcF6wscVw644sheTWt7FMi3Sh2/rGyBa6azFm7onZrIPv+c
VQIF8QMcPclXlMZeV95hWinM5JSoT3WEfBisue7yAtJbd7Pb3H2gQqDAiijcAKGu9ry5YoJAv4Pc
j5PrUMPb47omP0MgUBQAwrlYy9HDRLDzSXugkOhYOnXFqE/ad5ctqupVquJ4GDCcKGCa7kTqy96F
AhdRk7nnCACSR1x5+E6/feKcFq1mXLzwRFGbE1fgsS9TCO6OSupfSgX44F0DBGlDGhkWuYQ652Ua
ZiiU2mr8xefRv+gD5YcevNvvkHMKPW5nV+rPZtEYtqMVgm1+imNecVKVaqfwPjecxMqdDDcnrZlm
Triqw8aAIp2qODe1O6wmw6XI1AgkxXuA2r6CTJ1vDDdG0q8kjTVs6I/yqOHq6XMRNs+njvdWPhhT
bJ6z2afuo6l3dKLm0IYyn5wE/k2jqvZEtZSG4cFkJHwLphU+y46m09RdoPbPUDr4AmhS1iwRGwSc
lyU0WAWww45pcMCldSSonNwJvvPAYfHD4tAjdWGWUEaJgklu1LFbs6Q8z3H2YZfMPICsdVpJi57b
aYIO3uz2SAv3XeI/VW6lxGRym/YhyZT+rvVIYlHVFemOrLg3xvTlz2w9JwcVDdr3KDEnQEUEFv2J
LMvhGWT4yjLxMzr1u3SefqMo7nakuxiemilNO0wR9ctDzKqlCobReYlmcyVH3ylBurtpfXvD5C5L
Mq4VTncBN17vPywUaFWHUaSajQtYzKRgrOKa9N4KAVqW028ScDVGPlGd8bPyKxkRqKMTim4JSkaD
wAInsqAkhVudO2h1ZirUxfLnVOLj11HSzyDvY5UFuja+PoGhY5TP36bdlzIclfIYKtyhpqmUQiXe
aNfRPZN/gFoBKxcuflbB8KtOEF4mPzpOy2nUlIxRkLIqKnqlXY+NeXmyFKGHzeyIyEIf5sB1YdfN
AnIRS/H2w9YcEtDyj3spRRLMYduMks9DOPIe/TZ4RMagHw4y5jlocbl4l4ajN+QKsjnZzxwy0hoI
CTz1nNx8D38pXSPyVdY+sYYNwtLv6GWh3+j7qC8a+dKOaiVL/59/Ghbbk1iupnOZ7+EM4ohx1oSj
xAsuxQbQLTsLG+gjttGV75u9424iW0/tU4AkafafyDbp7WyulV8Kqd94k1a5nStM2e+Be/D6UhDi
KPzmeL2YXQCj4fmMOS/5iERPoPsvqPEtnNVx33ATMvAgezjmpFqX+r977ArgkW3WNHNs2Z3pgbI1
k28FbUUEpkM27otnp2LHJ7gmvjT8jhmfhKHdKB8PnDiUMSrPCLStiPD4cvFJgNnST+rZh1DcalyA
PYQ8+WV4meY1yTBbZWg4CelrRWoPUgCQo8/BT9upddHlh9ug82Eut9FL+a4ywxIpmAQnLg66mJRL
C2ar/1w0pn9JY7GyCnCuMi4PxX2JSCuTQS3sbVch3jaTCo0vFJnb57eGa+TR+tGfCZ0uXceJ2Usd
fXT5LjSb9yAASYgc+OB571/ymqTBXjVX5Ur49QAEamhDkhtnkpGSG8JKKBDHpPQOFSgOt83D3QJO
5L81Nk3JcY3rmbRT78hV7UgvpYk4LnitBcgs2PlrFTlN2tLYouHkuQQLoM3kir3JngqRqfMxyUAT
gX9pdr61lfYqbn8x+YoQ21h+4sv7HP3gu829/dMyJDWY+DO/I03aAUGUjJpfLfb+t4JMRSByOlBL
xYA63m/qNlN/QCyWOeCkwGjOdW/WyckPMxK0mSolsFdfjWcUlQ3EHs7Odr9YXHh88EhPK30QGTGc
SZ+wo+5te2fvSQhLuoaJIJPEeaqlsMFcPDe20CFQvsc93zmwTgWQdzTn9+J7UwsiJsJjO3MTwOKC
GCpM6u4+J7tWjlnr9IU+/2pWHQvPyeAVWs1WTVvyCL6mB7yqA3A6jx/Jb7muvSkFTuNTqaHIJLZq
rN6QlNVUEyw4u78XKc+15PqI+S1MwsQPZIeZqOPg6qnafMui7RmX9AGioxMfmzfcgDbMHcaRdDXW
JcfvBEFFAl6Nmg/l8kxrQLPi4ENdw+8GRU42xoiGcbNR6gAro/bNlD2fvK482ny0uRpJhiuwI0tY
4tgf42TgFbTvvCuK+nzZL048o/05eIV9xwXJEVjCLViJ6qqwet2lXGtRgf9S4uTMDW91f/zJ/vsD
yuBG5QlTtq2ywf7qewFEN8CIuT2RC5f++9ZwYo1nh6a1KX0EZzKIhPNX54fyvaPbduHQevhG3VIJ
R4P7bHwcxkNfqkc5ct04zhKZCgxN6ImrrGlld+gK6uBHfPxLEKROr7TldGXAi3HKAx4oBBslIQ30
Zy4UTtaD6WQwH5Di0+B1tocziIdvoTAnbEPWfkMr4LAp1zLffgQXTSj0YoWaHIyDN1LoNmWhqTu7
DfKHOQ+sUyA7HLn8FBuj/xXa5R2rdNlJVoRxQKkCiizimrq+RVzTFg4Rr3caCEhPlAr+SOPuNWVc
kvZVWwzmN+ZTa6y/O6/ZUBj1X2V8jDgBAq93+bo3LNnord2I8514evApRzsLznms+HpJCafXE1J9
fv9R6wOPq7ComqOR08VaOqsDIpGtasFhmRsOxvNK51oB5SvDMoIyIylz9+wnmN9TxPXo9IuG05/S
Ia8M6+XZBk26RPTqcLad7ueW8pxOBZxENf/2zC1jNTbQeuCSI7BJq2U+JsK7FPpYnkx8TFPwPwoj
0ARt0EOwWw7zMIpqNEYkv5yOTG+bnUi8bm6AgV9AbNTAlRRRqqn75Y/vyZMDaCPfzKjWyuuITmdK
U7+3eYR+UFmFUVPManEVAGl5HoDV86UtH+8qJ3/SixnVzEba2S1JOTTz3bvthsbXlGckykxAdATt
zSQPM/DhJm4Fo9rzjk9m1hsOHmH5E4dA5DcYdReYQWeRGlCF9cA/38kDzmj5pK0IsghB3TM8sF3S
Jov10Wzg+1cwueb+B99/GLhNh7+tdhKwld0Ai+Txv9RR3w+cXe3QOsLhU6DrGSzU2IxpexZQgEfN
sF2wbFTZ0gP6cqAPaSjSJ+WYrdIrku3eGZOGrVRMVA/XKXMOigeQhF6ZNzrV+tDwXpVKsp9CO5P4
taTrZn0EZtvhbbnzw0/jMOP2CBseZD7aYzjBwAJGUKP+R97sosKrJrgs1MfjMuWjKws8NNi3IOJV
iBtX9ahMtqUNq8CxLSH4CihOY9q0T5AAdF00OnHN44SisBhxqU5XBOEGIX+7JHOl45FB1OdmcMet
08aM2O121+8NAqda9OAEPAQiyOsJNnEzC4n3YhR9Ce75uxdSmrblF+5mbmcae4rWwH+V41SA1oeT
Y1GshEDBPw/Hz3yVOHAJqQZfaQJHNJD94aAKlD1HYQEu3hH55Nxe866my3RSw0NXp6t5//uPINV/
Dqp0djUCCMtBLj2RvwgGuo0oHKPG4rTq6vABZDpkd2/Xhi9ugiqB+4FGZj/9S15OofPX/1Y++ISR
hPqfiwURxGfh922G68HRlYHngC6QoV2WUDhOCGtnxKrnb4qojVTj7fw7wyjTbARWS+JNw887linY
y1/+WNPsfh/NzaXH2TqZLyAudLphgmvEGYlWHb6pmw8lRsqyVFkcDMvQzmguVflybUUWySu13Qzh
gqYoW7T6IkdFHzYWC4JD2PJsY+Ug2B1BxM9EbkT/6CPHCLf2r0TsCluolb6vAgXzNg9qqOh44WFW
38IOzyenxoJiKBzVPp63i7Xzdl2PrMjweL2fonFSuVZjdrxkdUiWRqrtSyltH5zvVI6BC/IRKOpT
hL7Pi2H1sf1V6wvMLWKbY7WVHyYeQ0ECbHYBZHOK6ho81KnEIm9TAT7QRHtK3cSsVX4iyRDmbmRN
PC3WMTiiHrRkKzV4AceuDhQLBoU3fpHmKPz2YauG5NWrW1TUojZPu1C47H8Tk7oQgdBfu2U2QgfA
LkifjqbMdPJIX0A1BAK3sB9dRqZpEhUTlcY4zbznGelcB0O3sr+amQVtUUpDL3HrU7dvg5lJJjQG
Z+kMvFOPtO0vGR9Z9AJY9uxvqVBJ9ypEPgWVzzIpnqfvvwt9XFg+E8cGrQ8BIfYVMI1uetB5BoSy
iZh8W5nNlnieFtXNj0u6lI+KdXlo5C1+ab6jHRVc9Q9UjbBoz3NtNuQN3nM/+nctuM4+NB1FX93A
cFuNMNYTCExP0zg+rKOnij5cLHTK4xPp8/dlXXP2wz3Wt7KJtqSgXd+03L1A66E9kACNIyWU6k9r
9UCN5UYY1xqOONiTZflqgvmBkA+dVghEDR/0y2M1XzaaC0HtymIeiEmsmvZ97mxwCYLx4PZOyHTd
vz+bWmK+jyA694RLXJWniLiZkS4RC+ROA/R1ecQqeUA32CFRr0ntW8IlAsu/qHbvri0I+a2SqvLb
g0ynzwynMO83R8xRJRusHDkcXH4Bi+IAO7vAxmiuuORpnTg5l52Sgqri0M61MUamzBxDgykp9Ok0
k+lpUzZmURrS34cuHdEk3ntR3II+58rG1xtPNg0OZrV/TASAfkZJvHC5+fP1mi2Wqolid4S8roMw
eXPKNXJHqerA8uo1zMTE9e7FxgRVc0eLlAXwdh8oHbXxVK6dNR6zBFIxKQPBXaGQdSgZme88LAHf
t1g3Jo6XXdmTwz/VjzrXblVvRQpREUnZnLE4jVCfBDr57G0itSyzbbt+MXzE9h/EHyxQZ/D6dx/o
+DP2xsYdH+fpsY5LfV+oDoR6atHQxvzjmpWoyOaepFTv0+nR78rHZRXXeIXWLn/J458OzhUQ01JK
tm+hTCJ5d8EaHHHb026ay/4qcvvsWgatDBAAyrKlnoAYXzF2AiTTWUkAhP+LILrGG1m8+cdbFumc
jyYS2BivyIbmaf49p5KMbwvfNYgheLgkbuX7gRDi+P7fAVNwVNzzDvPrQ86KsOl7JMkv7OOXZ8f8
/dg69MN9+mTE/EBtLVknKjvRfBdBPGMpCoeEgqvtdh/oXwnP5wUk42tJbG7cEH1Mzdao1B3tvgK6
PjynYQ1vBibdu1MIqd/OKQBBcoDJhQzyj/3bQwKIkl48LnNSGkCZCMlh85r9Q2WNk1rWms5270Ez
vgf9mQ32swiAAE83YfQPWZtCEiwqCf3+mPsNDh75vTdCwOzWSHy8c2Bw4h02FqUskxZSxUiT59WD
VHfa4uFIO2nqMfgd9CRSYW+JttHcYoIs5Pi99EVLtRNrJIhOmEM/ycgBGzcM4davRn5B0TEOmc5p
Sz6lVEDSiwZamHrBnImdD6x8sIBDfkKpTx1/4ekpc9wA4RnQ+OruHqaf18SOMUYIYYGeVSs/XHnV
F9wMA1tlYUynISWCRNGDGJdyfZKAymDsVkjZYLbTelvL5o05TKCuedOR92auEhl0aJO+iKw7M8nh
kWW5koYd5E/ZSjHfr42edemutLk2ku0Ru1rPchi7uaQbJPumDykT6uZIoSdE3a9yY4n77KZviCPh
5dTrYoa9oLFnWVqq+j7DcKioftmVBoudU0JlQ9V+XdOuSA9UZM65AAAJsXEnqOPkHTuNm/eg0wkd
4N9JpeO0QXRn/kl2I9D9oO4zRDkAW6V9jHPfHXEEDjW8hJG0oPoW0ivMwtT7V+uxcQ+ykCXZImEv
B0BCIi7G4E4ObXdHXFbXabkmz69wuKtUf8W4R7dS3jIrCR/V/DtexG2xo/z+zHUxfGpPlYKNXj1c
R/+y9WQAlzfdQccLA6lMXuyhIz2opHyKY5T88V1hw6keYOfEFx2h3Fy97ZK1omNG+EJ94q0C95N1
uaC9yNtIyMoFKffUGht0M1RcRdENFQEuVDKEU8xiM2EJQ7a6nMpBnNPTizfN9Ov0a/JGRn+UobQF
EcvnYI3i8CdjGPQ53QroO9eRblRMhrQV+waBIPYGcQBTJz6ZmUn63g8wNx3Xx7tRFrulGzsQLM7E
oRV+EG1SW066gE6IHqsUC59ptoK9vQh3pZyxNFBf3TBMr0enEt/5cUAga7YZhvwYLHE2UMePql9A
1CyEXMcuy+CHsVLkQLJNVjJoVPxohkr1dYGokse2QSx3Lqy+a0shhoaEDAXLOZuuPwiMHxi3ypct
T9UC5799B7oW1XLLtKXkCSCLtf294pL99Fo/cEoPm3DmBSJoyYue8zw4lmfMUZYluT5Gz8it/tV1
IJl1mdEpo1MCAATAdrTiPwNM8hkJVRHsiF6Q4qcoso42lScdc+3V3h2QgSlFcmTasZyySH8/Mdb0
KTXxr4AGivjGAgihvG7FFsIKpCum1x/EmvlhMhNWVe+oDIS2dT8v8e9FVEhB/HxlxDC+8YzseLhP
4WoNh3QOp0JwYOPUdJ4KfaIFNLUvl4TlJu9h7jRuVQtNvvEWHWQKJhZsLEk1fRgF76KfRTJX8O1g
q6IPYnKA3yeMK7PXg1s/Ci3+09hW1KePPGCbl3d51wg/wknRmnpDkMIPQO+Sn/MHAIormuhfoNJj
sMvnMG8dcnk7RZff1YUaEHh7tUgaZhxg/5buVYkKdQIsIgPBNcQXvC8DiVYV/SlUKmMvPE7Mafof
LZQfX/BF225XqMo2hdgcAdFREZjeusTAsk+rB4cNd5D8xLGYpYCgseWXGPKJ7RavH2Rqs6hYrAZh
/vur7TKHex5PJq5TMoCOI3bdPbeqAdyaDe5PtWMVAftUMxglEKAgayIway9FpZenoxLjbInlfu2/
V/YS798jd+uVXwuAJei/BJ8317TXBTCAwnJlRHWNtkqQMNDAMoSk8JVoh1n6VUoxv0Qtq1IZ/6EZ
YZKMm6lwA2eco8RvczVCuNVtkIKDBVeOkeLiqE+j9+AEFUkXuF4lEbxT3ukEa3bXw0ZU7mFyQ5vZ
y3mYaCT+mbiCXEojjXuqarv786hRgIoyfWdDy7vGcXn+48xse42AZT40mhkRsYo01TZyiAQR794u
7PBKA8PY1+hEVJ9+on/AcvUQSejeTtGjhOB9apFaoByBx0yACjHRis3PMNX8KSX3iviaEWnHHEuW
e0GTy5UZi8bht71KgbacWdw2DJExjQmNykQnIRi1nXKiLW5YEFySmXrNYlwiT2tW/VRptMd9bBrk
13nFh347nY61Z1WoX6eDFzCQPQZRKCAWuztEsfEUFqFj0/JdX7rhXh05BwLAUs6EdikOn3Mp88fG
mG+E06Xsmcxe7n9xOvI8va/PPiPIrabaaLVdwka4hTQkteMDYMbboY7NSoSx6FbQlwFAx226E/Vv
jiUikrY9PCzSLaClp+dVooy9xlxlKOV1TuheW1z7nPdFP/CgfVObJXg8H/t+gY6WJDL/lY8RkRkH
fw1FXFgb264Z4KiT/0ItWK9Df/HIRiSEIGNGAnAimYfLRVSnzAW6l0FNlTfmO34/KmKL2rdgSvOe
AHqRy+rMWCh+Pb35UK05geHfvWk9v0PeXpcdUUBbqTO5E+hhDELQaCqQO4Sf24dOKb+Do/sUop5a
LzUGEzwz1tdCh+ZUMD3Z5v9K0CxigUB3E8XjAiK3N9mqr5xogNMCVzHhkOQGZ32OA5GmmRe8qc3J
iKTw00Zx/+wzFjc+pEOAxACXK05YYBDtxjARhW46r6RUwTrQJHpn4EEraNRKIRwoHzMPef9iNhsd
QIrAX+2Nc10Se0ZDUFZaT5Rrl9OrAjJgENepfhAGhgqG1Ss2U6CcXHAsCSi/9uj8aT5BXhZn2fpc
FnRQKa06gw+DQyQ8wgSp3zOZf1pcpaNj3iXN1hdX6ViGbAI91BLvVuEjKT1idVPyPVgcwvVvY5NK
2KrlQK2kUraVZEt9D62RII39acJK6EWfn4i94OE2BBRqVzBL2vvVZQsTYXVGr36kwv/qjKVC+03M
Em8M8YVe7kYAPqlMLBYUzTh3lowRldIMhPiCIsGi
`protect end_protected
