`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AlIIr2bcQt5eY/wxjGFlAFVJWSzi93+Zi27zqOMo1YqCDQ1gUj38mwjC6XM55QlLNAScVZW273jV
X6kHYXTXyg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fdAyHKzPmAELJJGSTpCGrIhlftW6NURul+L7KHaWZ81Wi5r7CrwBYRssf6+vIHm2cDXkA/iH2HnZ
PGTaY/z1sWSLIQSxDZX8W6y1UiQtUQEnph+9sOVmYV0LrNMIYzyTofqHc2h9vNZAafYiQfVDJipg
W9VPq579SHpevheD2MA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LnWKV/dWXS96DVk0G6UiutiyAAfw8RxMejgH6QtoSAbK3FejF3snrtKdn3rsgOWeDhYAkFYA6XAI
cmW1l3hyB8Wi9P7FRd1DFPMhdF7vRIF4kw/33ZvoEuiJ4ngLuwHxwN/tY4pD1b1F5/pUUHdIW762
haBN/yKxh1PXuy2GHBRyk7wD2hUhguDSIFoJwYWjiDfKmbck1IQmrr2Wg5g07JVcdLUrLMxfvx5O
7kdl7q66Pfz3TQ3E8Wd3csKxo33az1CZPBEWsCF07iKTv074dKyA5khywK7wIkhpQeSPdJACcKqM
gKwoKGqWMgZxn0PjXvzw9SANxR8fSgSVI8sh1w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oP8Fh5FCJ6I1qIsFy/8MutqLA55Htt0VFGS5PDp/Epdl0fmIr6WHjGcVtleZhTxwEVytT5XuVL+V
/XN6ABr26QrOLq4yuREPEfMAllaMH8dEd3VZ9mKCsXaaeQhL9h9IgwvhcNQKYIVnA7+aalNq9D+e
KKVfCzXavx8P/gbKJrVVKtMQvgLacZy6cjiXSyWr7ITcJ974s7i99d5tCBCHG1XUBxxSq8FD4SBo
7RkYOf3+2yZT8gxlJ8ycx1JKksou6ZGLtQVHr21miPk3RV0MEktLi1/eLWv6lZweVD200bPCgdvj
mgzf9s2NoOtldo5nQjvVjUliFuYjiI66R4ICAA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f+ql+sEoZH+Jf3wGXM3X+UCWoPL4KHlT3TvjtbgIlbs+qW4DgNrI2ch/KFnOOFgqNVG66V6lSJe8
CgJ/sHGzVeuqWppQPzIRCBpfLe/04yHVOjJeuLx1duwYhek/bFeOZ76znR+FZLDImSe77ZlkWNrO
KgLCNXSkGzrly8KwRhE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lThX362nwJscYdxxG/MVse3OolwcldAzvGP3vb9JHJQC2zu625AkApJkljuq4hv+jyCvgdgSXxUA
aQ/O6YlMtyM0oUT0lfjDnl5qBjEcxlaEEFn/yuqP1qVoiPPKxAvRQv8o+od6AffANbG5VVvm9kxz
1ojDy1MxNv1hj2uEToa/S8bA3g4zN4wqFFVle1yc0awjYi1l1Qc0Lvcv/2SPBCMCiJfW+nuVtaeF
BdIU9Zm+dW3B/Q6Sot8hLfsE57l06WRLrSqaLKO9OFCmBUXiyXGT/MY6STfWOsd8vNjXT98Hbz5k
sSk5caLNq4hG0l4YG3ow8LIYUISZovYHZuWhBA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hd0vgBtYteHG7h7abWyZ8uuN39cmGpj5zg2wOAteo6OPyld/z5B6lFJqUgId0WuS37o4UjcoDd2a
EcphvKa81+U9OoVWFQxKXMQHisoQB857pupeG+DoUPGo+bUllCAcPbj2t9vwcJkpLpTxmeRLtj3L
lkmvbSSysWzH5LNORgJmWwAgQHeNDmpaO+EFab5j+YsnIECKYYKz13dVhUaPi+2aUF0TpI6xt5HL
y9n576lJ4geYPaRPZ23IxV3ZH7AhQ++uyJ5A6+aOgSIAgO5oaquDD7HZy+MYHOEKuUEIXj7KNcR4
YWTBmAp71qwjP/rhmEMv9V/u/5X31G4tgZjA5w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R7nN2+Zs1dKvW4vp0D63je5ydyoTDrsLefKhOSM1rJ0h4ZoJV4jZINArGMhvp/X+Bhsk//lGINdN
hyz2L9T+Rk3HVvf2szTdr1zRHBdrx9hYynAcAi2T4WOJH54HZZaavsnFg8hNyfHqdXHheQFZxb+s
fCWGdXboQJsbd2cMLQ6vX5CexdkF0Jl6OOnW2U/epbiCzIz8+qAPfWme0Ggqxl8/OoQrB+eDmG8L
j726bJSVFgCd/SNgrx7hATyyly0nwzCAAw1vOnoC6vGbi38tFkg9It9ejTJXZOWLwBmjEHFSx59O
t3G7gUg2T7Z+tu2G2CqNPJUw7Waek7sGAusriA==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I5HSCKt/WZTjyqd+HHhQ8suolwbhucn9B8G97gAgfO1MrekkoqVh6/74aGzPv7v5xutzlOBMzIFe
H8vYMVxUz4nQH3dYpc8HhGU98o4HXBE4/tg3fOZnoP1f01u/ztIyHfMuyEWpPOSgUfNZsjUNJiwv
djvLq7dSAm3l5C5bwZLCG0562hrGH9W1IPxJqb+ugTF9sQoVcYGZr6ob9ddC4CbI4ebtVFlM4ZeQ
RIvX822HYnrbwdFqnxMaJ9hNY5IJTvtoCqVKr71EWWWNRnH/OqYWcw92kqeuU0wJEbZGjV1dxQaA
MGezD4rrGAIsQLpKEEqEUxKArR8XTRaIiX1y5w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55552)
`protect data_block
BpmxSR3wAPCa8WWH/gXbKRtCzkZa3phi2OlcWcpbr1CN+StjYPVbq0/8aywQFjbTpypAjxjgvJiu
+cMsczULXii5+GKB5/dV1sgeKyBOVByndNam/frbxtLGcA3WlUF18Q3phJg2vi2pjfd2j0exLEie
EdHYEfKWrJ6NtESCr38rLjqDUAYHEMrYZ5I+2kcEta/vBkxw7/33ohVmLcMAR17X8Im2yEmbudhD
g59ga7zQlWBB9mCW0wvqE4qMPZ+T7aUG9DKeOnef6dcctLMlfWSUKEL4Yzp7PMZD2d867BF68BJH
5IRDQVZdHIuHm7llIdoE+DvY7iJkb4wgccpOvtdWqkW2tawi7FjaDqjbR1gbe1eyleYKFINGrYWS
Hx55k3t4rJ6OR52Q7iK3a5kML+hi3kML5ThQGArwL9nDJhDrrGs/gUtxAOvS3kYWiOPF8cwUfjJH
Uf67YSqGbkQyxd72YFuMT4mUL/tHVNHi+yF000BjijoWGfYu38A2z0lqM7a8ZIEIj8lRnrS1DLz3
2dpTXI+0V8UckrnjbvQycBBLlSVl01i8bVWRnqCVAQzphnrqDIYS9muazJiIrk4OC+C8ma9s/1yg
j1qQlKrxOgBpUT+KywfxWZ2WiBdRm994fahOStrwalHRcCbhrn08mmJxmAL6tutXr5RakPBBPKPx
F8zXEoG9d+G1JN1cqjO8YD2Ajq9zedGh1R8nHSFQwXbWJun9Vee2+pgya/rfm8/+Rk51kmSEp8mt
lQHzlhb2uBf8O/8FShtXJWe82sve4Cl5FpMpXIR3FiDlJrIeyLDL2HEm5wPHPUHlr2KUnWn9PgVE
ZQceOEvtAlDADPl79Jee5pKGtmE++9J2XHsChKNJgrvpQMsXk9tw9W+y1Ysky1kb3eUmMLzKeIWQ
a4TswvxBwMGeUgtiVb1YPpDkfhnfteaI4mEetvlZEgwE6AFzX73Oaj3qc/Avy5Ede8N+ftH2PtYj
m95hBdyWH8eH8CDqSOeS3xLEwRJknvX6Xs4M6asucuRE+zN7mqZ1oGbKi0EWZ6vJbHrqXljiR0ek
rfXt6z+SlApB6IVxwWMtSMWzN85HuvwaeC/orrosrHIijVPZ9gmA1Jqwo8YKwjA0brgsOhbfM3G0
GmwgxU0Pu7xgJM4Sfpym1a+RiVcn+dvnyIlLZ9UDd1rAxq6ZZ2teGzAwj1LMYA8vn2CgW0SErK1R
xqnL9WK8l5LL8cM/sirI+v4ZxASx1F9WlcZlJf1BtSZpJmV6bKvZIlnRXV+U9q4zm9//1vvx1ZBG
OH/ZODrn0yedzKinNbS78DQN6rugh5pfpxPmoRZlp+/W2lfms8Z7DMj6j7GOnrZqK5uPxLeln3LO
QWUGPz4qjDFf/fbdXu5xiPnPHdAxlHBkyFgyGF99EzeYTQek9lZsBpQggxxO7RudogYMw4VjEt2K
zI1mgjz1XKhMSQTD9iCGRsuYPDPvKj5sp4wSYZewIxT6D8Bdivdv1tMAJCzWJC6YUwynCABkA147
baPR5+mDEtc5APiXkrGj0lSd+/ZF11N17zHWoiVr/JWY/wRB5r6dPVjiv6CFaY1wH+YBw0pOtxdx
gWQzKxKviXFY5UmY1PM7cn2E91fDNY+kqK3q7hIaIfkW/SQITSsiV4SuGzsjHPo/AD/7ZGpgpSEt
rCEsEu66QHQTUIip3DU7MUblVFX6VlWXxDcvZLEKqslJHQgpissmz6WiF3YsKiMgQbF3OY5biub8
/QGKukFWcpCaG+TW6GbRrmZmZTWLUbvMdBYzcMjJXtJ8tt1OrZwLrs2wtm6w5ZqlrTsBta8MfROS
yZA5Lk1cb9OCmzgwiBwfekv1csVlBkctxTkArdUWcYJi5sHkeX+V3Fzkl6jL8JJvRoU+4RI7PXio
1VgSwf1clc0wcyIkx3etr3DAC/pZBlujDY73DOENU+8OJio9hix2tcryWNsXQfKmJKnGarYTpWTE
dYQ9Wnshk1oclQGoEof0lSOkG+uCsYx/3ZEE2uUVqkD5FeY5GImKCM3s0QliPitXCxpmK+++fyHx
QdyIg4xOdi0+LhrZuZl6snB7EycuKxCo+tTvaFhqk4c4fShuY7kkmV1TXqEmQlNMq315Vmj3RnJe
tylu6J+j49SmMy0zvbjJhPQSudF4iI4mz9Va8ZeWJ+27wQjL41rvVc9URtrFb6EAW5kR3NbYws/8
ILff85LE7XKiv3UP2y1uGK9aa4gFDXPoxosFR07Rut7RWXF7FtGRADaIii1/mb4P0o4oU024YCSn
N/rB0X3kgsInXLqH+e1bRFkTlL9o29MfEn4aayHhlZp6Xajs2p++SDh20iCe54T+eSCy6/KFZ/q1
svIWDGF5zDFK0OnrZ5/Pp8L+IcltdxaCRIaGzloeU8fwlmAeu1rikwyJLGwM/5wJhhc772jSllET
mPdNB8vtPYQYMI+/nPotsbkAHrt54jVu/3OgF8MXorc9GjxBmdgKDV8Z2QyYmWnEHYm8nn3yMdXp
pkevisNcpx362m9G+vajc/PjxUZFSDv3I7FEnZgBvTZqtXo2py15wEIUCJ+noEePW5pSWE8dbsV4
1EXrW88xTFfZiDyl6QWOvx7Y8/3NVh2L0XRfMYqiQ8Qi2PPB/3yWP3ixXvHF2gsjcfdNAhKk9TM1
o2hBGFbaB6FsVMmwlZ1ZY+viQz1YBdMG1AyWe1UUBV5ejKQVQ50BEub5F8hi2Q8Q48dvC3FrWmQb
1JpTq3vTZcEHMiiNwSSJrv8vxc1X+Zg+s+N5GcaIb/2TigiPvHUgLOyNdlwkXqc1BO/ReUDqRtvh
3/V10iARP+5wul8b7qDtX/CjXIkvKTqXXYgbU3i7ZxzvXJVaXIb1sQ1PAG1VsLiTcwN/0xl5dg7t
E1m0N3WNdEddTAJI9Xeupsm/Xj3O0vbQh9SxsetSV2KqJyQBOqU8FRvmZMImQPV+Me/K6JG1NbRu
VRbVbZRsSuLQ1ByWXlnNQ7Qsz48CyzQRnNJUqcTA0YqoeX3kNa3+ItFjrmMHVtUBerNMmyIkrWYs
MDZWHI2mDvCL9JiZmTmB7n6qX+lPEurwKfkbKmGTm90j7FaE0ckzZ099jZ9oQW9vW2TYR3WY2N39
S88IC0pCg9S2aHrHIYLvWRMlKB+LPD54zCNrcBoCqDLO7qS1HWcOAF5M99V66LVHLKM3ltiMeAxv
LYViVg2E0s6hNdo30AlqJHWnDrP7ozsx2emVTKlE8CXZmGYq7zMzPBE3r7rIbLjDQnKYGKn37PF1
Jo4j3JJkd1cb1AuXjmLsMIKQi4YFFYR2zEj82xJYyPivaUnG1CMYwnot6wLKuvHBg9urSOCmQJwp
LM1PfV+XV0hETRyyklf1zhbncRv0BBjJeYsCbnNQSLN4JrAU1KGbopOTS4fOFMy1I8HJKJq/bKZI
x/RNKnWx4CIEvpMQaSc3t5Wkg1EHuDdgCazKuL/dYSDjuJqhWNjS801oogGVUsC0LNaO00Sz1IEt
wEZzK6SSbbeiBc9BrqNi0vibuvheFZLmXXffVi1x4PIanVJNGspSpsw334J0WXacZCmvbGQQww3F
jY6aG/awCBM07/LF1swUGSi+h1tTSCDQb4QwtxSfe6TUeKh/4A5a1GYKYDtbYgyeCFhpPDQSjPSF
p5B+0c3Pe6VCwTgj9guXiJljvi1MCNhmZ+68X29PSDgl7BMQlTPQIgsrW3Llbeu7uN0FVJmUw4de
gPCoxqvXspfCmdZANmCeIGSexgx5ObNZiRnpEr7oolJZRo9XujsROUxHjF6/mA1by+TEw25i7qDI
erbTETRg6N7n8jAQwctpiI9tiqYVt6KdhwFp40PxiVbKb/SDCySyZWqiSe7Icm6lZ4LVVCEBDr/W
q+a7CO+DKfr1qZtvChPVfpFyrsTxt7Wa5LozOYP7aZCbMAL07snh/UjG5wANMLz18J0t915JQy0j
70sJ27Wxy+IYx2EjnOnEHtARuFxv016nfHlegRjofwOkXW1X4DE4Us80Ee1d4YkNKm/n3P03U1sY
uthE9/5Fy00TEcGF8uIgTniawnEOW0EqcIyqG6B2ivQPT4/YpDFgT8Lze9j8wocnmPgCE6w5PIpv
F0+tGZ5qNrJq7hP7kLpKMiP22MPf/Q8pZnUV83zC3aQKQSeXuKHGaGhL3haw0CK79+5BYrgrqDCW
rPY4QrNF913HJvnC2vhOlFf91J/DO1WqjU9wXWZc9GJrruSeGYLZjDWjgkxalhx4unA8t0TZemrq
P8cxzvUue0hxHH3e2X1s9FbbfaEpA/yg0bzF8w4JUEZPASdJxou9DOEa8FP3Yp0TYOE9+HBg/vMx
CNsQR79g6pytZUMU9ho24Dzy+JGtKJGYlfFsorswLU/2r+deflE4eswv5LwUTR8t8bjSN11W+2Tk
JsApNDnv/i0MI2ZEr5EmXD3trVraJOMaBpeOdP40TxxgrJXKV0dSKrPeUve5wxsESl+7ZS1L7etK
sbBpOQoaqT0Rh7d7sr6KWKeGIpmS6KWA43LFZceKZLA7nY4DgQDuVFEbZtXlb1iorD2sDjMR5swA
EdVIER/WHTstjHLnJ2ers4gOTVCPb6SVM3KKVJq18dTSsVTlGGlI37Qg61xKwJhG5Iy0oMCMmoCn
xLVbJp5FfLp2S1SFZipQjypGTX9fwGvpmoupdtwmOfFHvCXltNC+9eJe64BWjLzeA/SkqUPrvFbw
JiZy4zBjLcqDZy9DVo9EvtSi8TMlmqfbgtzDbPy0ZqAKIEw267uqV3xriM1YQa1tTjZe6sPPVL5C
uwk4Wpljf9j8d0TGPSi6B+UpPgFROxmcQXmwGuRFdhDRLAZtCmWmljNpspVfvsyS2dTHO1wXr1+4
+n1FRnJNaClN01MlzWUTZ47cZWm91FKXT5Dp446z8OOas34HxS2YF+E8FPORNmU/J/AnRRKQdqBx
KZCAWfNiYVimYZXwNT1znQ0o3oUGLNmrMD0a8NsjZNnRmL34kXOfm24LCkTwjkRI/2zkM75MjJtx
FnaKafd6vB/1EajmXYpv4sumsEsE1xXatvkY27z6Urn3YtLCfEZDcofGUj+hVHQe0/ARR+NyHAb7
y03maZGkuD+ODN1bp+P25+OHIpMkacZNXJXk6Qj8yPS9Wqlc6h/FL+ieJSeh6ZjcdeGdu34+fUNj
2hEBk43PVMfUh6Tzy/RhXGlhcwNO16Cr/sX76VEtCHB3dNNC3NxROZXmRQ3AdjZNch2tb5tavCps
TNgmbgLc6zFIg+wjIXhooB6z5cMz6I3Kycxxg+8wkSNzn1Xh6H3m+56av+ry51Yh2szrGxiCG3Yp
VPJfJG6FeZ93fFMcPvYCTW0uwPR5TYynL6ixR81jydbT4jQKDGREfMwIh4XYwJoOY3Q1a1Q4ync3
jBuUby5eVayOyZhx6FGV+SqHqk7fC+TotbRLg3QV1ufiOrKd/7S6GuPyifOced5AYLGv3UdaOD3D
8bt1DavB7x4cRSHwzzVWyfAlTqlXTId0vWGvA9hjrRc80r37Y9pwTGF8hBlArAB8Oyb0nA051sOJ
VWUeOs/r0l74QOjBwZiXlHAOWFgZV3H8wOabZsvnTl1OHPXtWn4UV156Y8AdQm08SVbGQ0EzkoV8
VYaBByKNHMxpdE3ch26nrHa+C6lDdgmt08O0w3+jae+vNXzmcLNLcFw5RMAdBwV8tukQ+1oL4hSz
D7VXf1dhSR3EDWz5swjZYQUGJbT2ss35Wh49Ja8MEPRVMpZVppJ+GyZRx3PihuBKwalo4XYpQsHN
9r95IK0lOrk0nvB414K+FmNs9inlJGkwo0aF1tIkaStyZaXVlhtgUFZzmaqEilb9EKBDkxOaNtR6
N0E3RxjMfGAMa6P6GUkgEYrLXOljP+5OKR6s12Ui1w8mFbDCKBB+XhTNKwNMhpJnksMqQOZG4zTI
DGaZYNNFHui0C7UY98YroUFGVRhScWp3VtV6dE6Agj7rzqv3ttQnXQkpyPwPDb1BGQwaUX3Ww6rK
YrbxkC3EbY5Gpb6c3/W2hTCf8CnPBSWofi6tXvG3NUNrHwfBuBEqHDlsxmNLXTvnZ5ubme58x0Jy
RgkGg6KIpIvPs557BxMvJnuiuIiTfAkf1MLJ0UaNvvCWZVfOlQwu4eMQCMks+75xF/P0vbrAPhtm
kupaetiHiTBqGdLMoNmjAoPW1pUGEs4vPUIleJLcLbpEw1HR51l88Q/sL40puLjm1xO814V+3Pvl
h6GCLLoP95M9eHWNvT9pKqAUj3RXE7VRDLof8UfZgEJokeC/uLWSzwWZYm9JTkMZeXPT7ahZBE3S
vUOVQP/d8F3mVeAa0wLaE9UF1YNk79M2vFIzmQ5irPY0XOuaabmfADzIhQjypA5ZONq68N1p5v+B
Od/KF/Eeli3TboIKOtdbuZBWR2Wq/boWvJefi+PDOuit2BusArz/an5TfXwyGGq0XsgekyPx+El6
EXHBkitdXSr7AXerL3CMf/SGRT3rknlpypTmhbaApVU+PbGwu//yWHIge3GHlpS66zSO6q6oSyMU
vDTnPE8fZ8+1TIdhQXY+J0Hm4rwGTYL1TubAtPFjv8GRMjSihWWgJem3z1cBWDxf6PRt8x8vCurc
+gyAJGeQG5WpmPiE1OCD2xdhHXvnSrvxopDozNqqIGCaHxDf127y0IYqbAw31XH7B8nR61hoiYY/
NK1pU+TSkxy7+5etvm5gtxk6nopSyXZpfQYj1kvHWQ9Zk+FwvYsmiGVDsU7wrMzmDLGCRn4biHS3
hY2EINB2t6SRHv412ZYHVkIUdwNJh1pcEqcnMrs14iljg+6yUuImwghbHdhPxnvlfx19kDXi9lQm
nhUXOOQ/qWaWxyJ0rTnTdcgut2lLGHcPT6eP4wHmlMojrSpL24kfbPgzEGsBG5bWieo97emwKLlS
M5jMcFxEEaLHt+fd9q2JaNsaTSpO9OCBqO5BPOTslFOu1ygVHR7z52z1eiloHI6Xzu3mz2JxdbtB
qw2skaFDm/BT2QeB8IhJZludK4WN/CzVCGkU7QoIwzyOd2zcNIsqpQIDGhBQ9LXgL49vrLPoV2H9
LrM5hzmpuRyx2R9yy4kr4SUgvkUkR8mn1G8UdE6G/EO5wZgk8sMPFHMyUINBDwS+MDTA1jhMlYrK
nHBhSGoRw8QbuzlbgWrf76OoEjQamiwjnCWg/TnetpFpBft7fwPcTvTp+WRC/1szcINUxQmRHmyq
tAX2VqKi8on7b+wGoLtYMYd6jFOrSWFE7dYKogybPy/N9X9xYHiNfN04iSHVz+bGiUlepnp6z3oP
epyVvvLuAzzyt+2FfxdraGvCuZQFylYPhgszvaY2mTTuyQBj4nqnBGNuCZF9+2x+NETKsNrNc7m4
SzipBbLtbV3ipb37ay/0w/i96wT42cfi0y92BoacPqDsLVKHCZHq6HGanL4a/mdMU5ElUcuIZG3d
XIjSz7EGCPSTUQh/yCmRjHvc5z1DTxUs+9wRJy26c2MM3npvjochWZYi+0EX6nQV0CJq8kBNEwAl
yDO5PMUTYMW5IGhqyiJ1yvLEKSqf5syAM0jwPUCXDRtsC+pSfR7wPBJlwYQKH8PpK/nRntN8/RQs
pckdV/daXD73cwnkeW+Tddb8rF3e9RA6EXYGQKjVpW9zpttZe5t7wF3i6gySIOzeWmGSKzraU3LF
nSkj/Elb8v7dZnAnC4xnWzBnSI1YGtrow8eZrZDiBxa4sJL5gpiou1fTcQXI713fu8EU11grkE4U
9TWhMbpXRks0ls2GQcd8TF3tA1aPW12yxP3pNT1CVjoGGvPXHpAti5nFXAJZiGgc1T20nl/UAMxo
22d+AUGrx2rWELrAUyocWW8jkMJuuimtcttj/ouyafZ1U1jDi6C6O1EDjbAQ46380K0ai51NNoEi
GXnc+C3o7Gs5iey11/de1CwYjRDIqSDt1rCfsIG9Gkp6VBhvupnvPW2sHQ35J961d1HMLEX7TwDU
JDLRf1eCx4AaZqsnKk0Cc5QU+gIosltlr0x54s+fN2FIuVgXLDimdGBYnEH90EEqdrHb68TydBrh
zzPogICfZAVgjUzQLdvREvbFWrr4DkuT5sX6cdE2QleyzQmdupLrKhgfQeWYTlMB7xbFTvy5ReSV
m2wslPpFofoiVeQLOXEUiyUp7S+fSpip9c2/8uCz3KHzAg+O/3aBpAO9yXJnahk2oHsY4UxTXoWt
fc32OwrrtauUex3wp7AKoS22eZXne72ZFxaxrcQV8IRKH5DOmja/LHray5qQCcP5MCD5MW+9rwbF
T0AkaBOgh6j2YpeIwmW8Q2nDhwuA8HMc99yyUYsWwLbOggwT9br3eMIcvYIMdT0MSi4lTK1Q+49T
5eDstjJf9AenjiiwgQkrsr6BhhFhVrkSJ4ifXK09QsX6grXcI422swtYnEK/pXr2zKtWNTOY79OX
Wjpbt7bjsIgdQddL/0M9eh8BVDsV1dcbU65CRzuZHY/iGcI8ZSU8FUy6jpVbKF9uicCVR7IJNIgW
CQQ+0UsgnS4qKCaZmlxhOgLkp6mzA7/reUpcY7EgngYuGHsnYDGelk3brjiEhztmpY4yoSuxSyjg
AZbYfuXPoINBCCg6k4R6nbETnzob7SWuhny5gMAeUlujJlrRmx6Y+Cr6qpvus7rhw6I4Kc4utqcE
TAev4c3jpXGShmXFe80RqdAO42bldWGCD91SnK4b1dAIHWveC5MsACzZhkabbP7fY5EqMVla5POj
mgH3JBcOTYC1+XteXWLxt3emHjTaW2xMJvDiRnoA5nO//tn9uKBN9c9XqzlnBj/g7wTX65+4fMeW
J4kDUKNyVZYbvikTkVpfuc47VhmPzRrJOXr4Y45CgI/vjZLthd84KuATiqXV9D6ilisGoZwE2VOZ
M/s/eiIeOwNDMrgjblHMZLNBzGWi37XAxxHv7N6FyACUbHbWXEjyVyItww0qL/y3sm204kFcggqu
lI9UYlif4VCKeQ6t8GNqajlCGblI2ttri+D8Uf3hgiQJ2tFoUQXJowMJznp49rkdabzWV1ooWTng
tG4xkm7XGBisEDtfUav3NRXDzImMqX2sxBZ3bdfEID1yLCD8VCVixBEUnfV9RlBageQjkqW3u6Tg
Rn9Tu0bDtZinYK4Pb+sKYMZV2cqQKb/i7W/6wpudatJDJGSfymBXkgRuIf4VDZJA140jMmlbK1kb
ICmxc5Tapy08WeOxXj8yBT9cNEpCNTy2i6q2NXOVSHk0mNElP8TEpz42GsLB6wfWXWe87dGx3ILu
ETClU2S61vaHhCu6AecNRf4H1NGADbh93V4IwcXYMBuw15x2TGgfgrmiYmyTDq0VRdQc4zDrdRX+
0/JA3Hq5tuAdRzOGYqhKIujfQMP7Nc529KRZz5BHIjnH2prNr7cRWj8T4gEkN0UoEjD67Ca/mYg/
WK0sUd1tM3Dyjdt/afgvLNVFDRdZFqwTTKEoc6Syz8b2VNALbWFi7PthSYWgtFPJ6uSdh1WVz7ZC
+6Pz4WZPUnc8wcgmkjbhMDqf1xHhJi3dEdjLovMK8xg8GKvGSxRjGyxLSqPcEjQJT2SSNyuBVZZg
2tM2JgNOTgHE4gWfQamSLpooCmUHqM7lF5apVSwjs7d1EOBXdFpB44TCGn6w6drmUxxyPhxUePG/
2ISsDK2DRItpsIxykff2L14hRvqHRRMkH6A7zZ6BsnM4JCQU4JAw91nyZG5zwBiYewsRfLCbzUIA
Jfpjhtwi5HRJByK9dhYv4VoZjxlEu72bZLU+JuQtx+bXUfakY5LNTTskVaEbq/JgaZzp8AXrk5M0
w2MWb32nCBPlSGNJgGP2FJw7v4lC4zUHtyOIBWno7mSIgu0BS6Bnfqvwp1TO1Q1oszkoyO7gLtHv
0fY3B8gPsMfDBfB9i+hQYXc7t+xDX4hTbIu8Uy/uLNv/0eajOx8omgnhPhJhzT66B7sUVJYta6Hi
rKqnlqRjowcYdgYz92KIKOCKzJpNOaxNwdahJhBXN7ZVBdZFHnKhln5LP5Wcokdwy1jC/roIyBZU
8SAX9KuwdqsVADeshrSWWxEMAR242yO2sKIxJi7bsyruxvsT/2Ol4iKI0Xct9arx/HcP+eEx+lMs
IYruwNGXV51EFGbD4zBBeFL7Euze4nsPtIVyDVzeUV/3MQ/bL0yyjieGvzoy/vF5FIENboEwJGXu
jj8NCP4Opw0SytsamKOCuCVsDhJ61cp9Nbh6WrTOWHaxx8ndv5P7GQI1miBDlylapL8IF+FOPWlg
X0fujfV6Rj9HUr0dFz/uNJJjkCPNKyZZyxmq930kVEdjpZAr7PALcGAg+0GdbmGPtRoAK91T7dTK
KDYISeF3Uhi1Q3KBC/XFfIJZXhS6taoqa3xb3fmelB0c/zFa2KvZ4YpRz7I4PgqR1uj5TOnq/HNQ
rDC85h3MUAtmcTImpan00bUV/Jd/3fD/G4kV+mhwtJvXEKUcXIwPkSDzkP8ixTG51JKmrtMg+/rL
wrMfTEMsjitvGbaps5rfnTU18KCmAZfl4UVuDQD9g3xGGbS88UaCagmHJ+L3en/1uemu6BVORWMd
SHv6QmOPhTdN9QZ84mk1PtnSAYFwUy2oyJavKWzs03ImVy7PBJK+PbGRV3gzZ3z2nTV1X8NshJwP
1+3WS3wjcczk3BBEg03ghi9OIS5WjXFmm3qgoZKDjRkF1K6bZ7HwVRoaYwV2imdvEIOnBapwd9e8
9IaudEiNPWCCKdxNk9Z3MB1MykgohKgNYu6XI+Rad+6JnzBFdHD+30ci68NDFN3HEUZoSkuy8V1x
HZ0yNW5+juGVadZQXopbwh2pk3+jIawzVyLxkiJrH+GtfI5fO+ExMLWTTdbNHs/F+P0BChuhftQ+
VXGWw6C37p+z0u1sX2qBxb8ju5tZDYrxwEIep7BZiaJ6D+e5c2/pDy0LHL0Zf5QTPTtZH6LwaWJs
5qgiPGS0MDbv0kxrohPb56dTCAxpqF5drBc6n+Zcy9Nj+Ueoizx79AI6p/AXa2fwLF2RbGF9Y2YB
wW9aNNPrOTN1QdgAo/vMAaIg2w/xn4KwRxheAimO6JN+Q6Un18325M3J3/TvYn4MI1sfsHPnulaX
g5/0g1D2BEJ35SzXSARaMlLM3+ibtv14X8l8Cg39jNDjI3je/28qNWvbv8KME1LgYGPYtDbXxbtj
EdO5/QPgsEW6O9pTE0oyfSVLHtu4M42YH+lgE8S1MD3g4ELe/5thO9gJ/YW9Ke+LwBETbSyHV8kB
1hz7pYmcwTTlc4w44p+raRswQ8ri+6P0aI8x2yBzz29Yuba/kiwYjJaBaOIk/kFxexWvwbXtIzff
aCIUBDhv4ZO7V6zgCocA9DMOjKQSY/kwHntYqQ19JhkB4ESoqG2qk1/L9QgP9OQc7Cas1Iqujd9+
5q5BTshWzwdUMZL8fqDu2GIFr6s0XeqFXkjRmownQGCsvZbU0/XAg6ObqRSygXD8bjFm/+KFrI2A
XzfKLMFb5Us5p88UN2axZV72lxQg3xvI9IIppW3bfL2XwIdvtnb0kSxxbeHHy3X6D/g0/2ckO9uf
JVDt89dxl79Tz6uvBS/J2bvYu0xn0FTxXOYsFKPoqjkrghwpPbXGS8ALVX2LPMv5CwXfHyVsxUps
ZZnZXa7+OB0Qrj1/ezKRRHmEzmPlv/HpXCHECWEDBarPMlOeeG/hzdBl7UGRUw23N+/nFbSQNWqO
NLqMIK2Kh5Y8YnMhMRi3cock+JOL4JT492Do+hoNyPPatA6lWIlY/Ju2YUqHFeAG8T8HK7zxHacW
YBWqqMHEQymv44s3HNF8wfAHl7Lro5k0B70m/LMbhWe1JVZjfVeRcdRhxbCf5dZoDcx5D62TWK/2
JQ3JXYr/eSGZC1QFOx6VOjzzbQ7vId2y/CnyjANNSNLe7NaNaNSKzLYSXO8qqs0ai4smbp5/HV0o
EHkI3CS2LQo4E/lEyTXTou+IrHV5SFwE+noAgxzk2Chv5kRJzycO7+Vq3KuRduhEmlcdxN/8BfzR
Bet3X2gC1uWzbxhb1eoSwrgqQdev76HeEZA6noCUHRsF+D6sXSEd2poW+foys3vzwH6Cv2+Tp+/5
x8kGECTTCLVSdIAVHF7zXTYzk8cSpozw1sb/Bk/G3LzYGrg5WoO/NC+07i1FHoORmC8jFopOgjOF
Rpubi5QJFzCW8+GrKvCk5R2AZIEkq0bq7MLBp64q8CMqF5WbcyvmxkofTOei8dWw0eoMXlpUVyiE
udaPLXV8rCUx74+Xrw7q356dbVwNkrk7oNTlx+UsYJnpANwV4ombuNTrYfdX9k/SD93kgNTLov0F
tMX5cfQkQRHUq5Ayp+njw8xH8D/aM7eRdtAlreLdHKj0fnn2Ws71NspUAtHmrm5qRgIOSU1OOZjV
41aCx7391FVibBm2FzStVcuUmZGkXMy8X8j/aUC6Os9I2182/shq8o29Eq9pePQuXwq4E/zVtzCV
RijUNqWPbWeMcpQ5VcldHGFw+wp0yDHzlCBGU5iqTQVTZXy++0X1HF/66nAjf7AnZGUumA7mJ+ML
dye3ZzNYza02kk1TKCoWBT7XKvbEn4P+2zuloWgiCGcjMzZqR6KVvwAuxmdxCFpey8cAFRnA0kXt
EB3bdgSn8vYFne8q0tVuNL3DoWDVmoe/dZHUUjB2ncnB3qnogzZuVJpGAkkXOmmVVamddiwP18UP
vN/mMLcY6bJc0K9QQPqp0cVpwBllmAycX7io2m1Pu/JBrv3hlmbfTYjVDCNJsN+VDOk354hgk15A
3Dbdkf99OMQMMusdfRxj01tvZYL9286pkUfGgsH+9FGw1xMnQCjDygTI6NX2Cs1ZpjjPbyy3/ExR
+qt/vrMsj+YUh9sEO9luCINnqyeXjPMuYIJIVnpvIOkKE2gMg8PLoWmvKBV1oGrOuJEAGW1Rd3j0
2qSKwHg6PilEkGpbxjF1u5a0HwBHzcQxtvF85LN1K0ms9z/rtOzb0hmaLEdnTdERt8jdNdKYOgMg
fTirMVQdEQ2JrDrHvl5d7ydoWCNnBmIxtqw4IFg2O8kPSHOgu8Cna5xCWfCUr59dUlZVf6jAJ+d5
txRalZ0tO5Ue21sINggD6ZnQkLUjy5BVninkUmQTEnjH9kjTW+2AobnQ0kUDopeIeu94fprLiJ8b
A3KaCRp6yLa5fWvEvxEDmbC5oDWo2RP6KnBKB/3znYDn4o+Df/5IZCOAVUYDbwjXukw49gopVGqP
OAIEGW8k/JiLf9Nx9a/eFDMPoE03/rwvff2JBZG4hjj7R7wMy5/030zIbXGvwgZRL+0z0zYvSKEi
y0A0JlFt1yUA9D5GUpRykvfJN18n20UTiP2Vs/ogIGrvbgUmNQeJGxMSEAGt8Qd5QgnFKeUISK7d
mmtzhb8Rd7dvG0fT8EulD2b0TbE2QsJ2WOYg+rn3F3nUS3pWa5yP1V/VfoIOGK1qGVyLDGbiVVRo
iaImhNFWyA1gPJAhEReHvSfLQeM05oHhMF/Hgf5UnWSB+bXx+Xrb2dWJh97Sz04iirkmiuAOU16c
LH+FmFS+rB0cZK2miUO9ae9iMD0DYBEyR4VnN+joIiAZVJs5U8KE3vXMxDx+nsuGZ31EjkKQhL2u
9qdvDArAPJs2JfwZ6k7tg89lg2RHQWYF4C8YCmCiQgvPniFh1kugzupW/J12eritWTRBq8WymGVm
5cGzbaPfrptDbW845957pQzGg5OD0KNWbhuMp2oHtPSXOEenmOw2W49+imnnqv0wi76hudnIdeBF
8GVAFbXiUJs7c2AzP++et1GhSUq89zbizI7665EB0ZIIijOtTotSKeq5a5ggN/r03fAIVRcMjE7i
bJkVODBmxaEQ6eADASSgUOaUrmWPwqHhev2fA38XTiFZHGHUggb0NchPPYi6FCjT83QLseXagFnt
6kB1I3DKjU2KDSOAjGmwdpF+v/RmpnQsYB+cDSXWB1uGHwhf1zuX/1lW9nhcBuhN6PlDaVQCAz/O
6sYAl4Dl4Ksmwk6p1Elkn3oeam/0hVgqDrvoL7eSwSoMs62PENYzdz1BOdNd6DQdEwU2c6FjtAmR
ayDtQphT+481KKBtNNl4h02HBh+u9BnXzkZPTkfurIPwxdgG/cMKS0dGTPnrNjBtf7MiGe6C8Jir
dcUT9Y+DNvX7FjRDeF3JrH923yi10/m2GW8POhIWQRiinQheSh2ghuq8bWCKvj+y9bJN1sflorP8
p5bnJlZf1sS4c2GlCDm6JIoYTYhLDiXPJ52NnOss0zcgeuAHWvM80z3EtQR5DPj/z1asWp3fdWi1
mvbOLTBhkaLpnb9bgQD56VAMdby6HdUOBzwoYF15IUCGRFEsQ5zVkBwLPpSr1Gmw3Box7guK8CxY
qUlc2QPKEue8Q5CnIGYTxqsvg1ezrB/ZmYvyf7kaBmGPU0//tS+TO2sd6Ivx8PgPvdJ//RTiAspp
VITh7qlR5sLezutmQf3QTd1BUaC3+YgJfJEJFxmcaeXkvkdMAwBFhR+MYicsXIvAzT006uOzNeJV
OTuew3b5s4/BfHx002Z40kbuvoprJ6/1RxuIncq+Bz8ZZoABpxAClg6iOUxEo/bPLoeyU+buN8+e
1ffd1bXFPdHnwtj+BawItt375WmaOilgrbShtQQ6W5YA75BNQdVylELtiLSGCbx/lIZi7wLDHyto
JwAXRHd2yiUMo8B9l+lZujExxToSyRg1JxqQ0JLSBDzb4+T2sd+5A4IJTTvbGuYa+4x5Q/Kdt9Fp
0PN7wnhJqqqhknMsnty6mBLnP1fRMxxzv7daq/q95KMMJDQ+Jno+hYzh80IquRT34Jc/qrWymwjO
vApYcCoTrY5yTKWIZ7pbYyQBXtnphk/4WovIVAhjCO49T7vREjVLzn9H4pGfGip1XHE1cPFJw8rr
Jt2GJch12Xv8QurbQl+g+Vhju4Qow6eaLIy6HidCDamndgtrf0qGDOg2rsxnXZJEkSk2FV9kNBa7
siBXYSBOvescQZSv0H6ypfyFSm6BLUntkRXfkjS6MahJ4eW6bv75hMMzW8TzRHOY1rA9AF0f5q8K
hU4zXzH7oLmkoZuxrN0W1kdMsNawAbzYQs0XPK1lI+FECollypGiqZE309Liw0WRwGBTRhQT/gqI
TaxU95VJCUJ2fFs6zhRiLXtJXqMVovw+qC1KJwAmYz3Gcowjqsg4kj3PK7XVwY4vXO7O6/q0N4PO
C8h6ixp7NfH+/g54uRSNlC/t4iSh0wTtgoDBH27lK+UIKqeZA+Ld6MGj8gTM/XU4FiMgvri1SBxh
JNJ8bie9mrlkgni/ZS6H1Axi7z/oJNr52GiOkmCZG2dPBDYoQU+oZWKjftcQsGriPTENyFXVa/nk
HZOJ1JbmPRbFGYilVrBlq5PczpQ697NRnNRh3biqXnbgFBpWeTUL+/kI2okTyi2Q+G4f9lv4rdEF
MPW7vkHZc18euCVeQg5Wcuucmqo6oDYwMcGWaGyz9oTxQwkkss0tezvVrQivfq9waLB0WAIeQa5M
6LY22m6L2J2+xcZo4gZKkl/h0ConijB0UytLxeIuSwb3IOm/4FTXLdE2ejcGWiwJZ/RNA3DWTtlK
qwqA/GkkZgnHpPIMwokRs1uaB0JPrqlrPKcOoUjXCmYb+deu3KANFSzPYy85eYibvCqwf6lSaGyY
ibSS5fS7nuYPowdKno23uER8cgdCBzaB9ynK3b1+7fYlX+sIxWQLA0OPlVo0MlKMmOK9/y5DlCnw
G/zCttr37mcomwHHl6ttqWB7IUNKFsJ3HMHRR0PWFSpotVH961d5KKPMvaAqSrg0ilPehtxS8LMK
ZCjzA/NoDSSutYXfnI8wDe9Syx1Ub2CwQSv9ts7q2CL/qkHhiyl0PHEihS9tKXQIu7Lvzx8NzR+P
P7lxc1y1sothr/B2ZEXY/XfX+RbZUagGKvSxVcgfa7iV4rn3Hi//0HFwuLMmjI6cpt9zzuwF8czs
MnBU3nrYxWIwOFJ7v7kngmfgiztDxWkYSa/3XAVMdOMdMfTqAukGi/1Of28UBWMHs1mkrM8QMwK3
G4fayEhk6IXZ5Tj6jSh79CSgHFo0Is9DnLC/SrjnxneBax6Pk8QOgeRgBLaG9M+MqAc1diDGvWcQ
7nZqMZlxgYvP7tOEouWE9oL6+c+oz9BbWuLsUbnSWE/O3W3vMUAD4hDxw1px7gEr7M7JwbU3uhNv
/vv42Z+ZXSvuAK6iMT0dhXBhXQs7iiyX8QXjgeuh1Hc+5cdCamiABg62XT1uaflyXDLuRui+aeOv
jCKUn75ixgCWXvG8IL9YkQiMCMcMrKUCZcAlqz7PxuQhzPFpq1tw866s1bc9CMMuGxwMSIIJbzfp
k9I56+5DNx1o4tzAuRS6xPy4OXEOtYBokNH1QB2TmG3orpPCtb8L6memsLFr1PKpAB24OuKGtGGz
jn+/USQTTE17bxCFyq3iK/ja3dy7Z1FxG5NzVI/ZnoDcBZ5PQa14T2I2YW4UNVKtT0EoYKmBvPcB
R47qu3SeZjqoUTyrJy3ojW/Wi0JGnZrqmjWBRiIJAS61dIConW8maUrzyvgYmE6Mkc5vDn2gPL5G
tG02wIp7USJlALw8All/Ch1FKvEl0OYU+1JX81FN41N+HDr5CKwMx+g0O5g21Xm3oTgqcEDzeEc2
9chEnqRKoTcSVGrQXkTNAKFlBc8FEMjHasCuU5azvLaOIZkww1sBJclZfxVk1gwZ4Su2swjev6pF
IhIrAp1NL4sPaRP5iz9X/5oKhk+Mk7rDxm5rO+FWFQu3EXbts5f3QMsKSEvpl8YaWUogcdkoNn2f
u+s3GQJ5zef/JPbjMimYElTGzRRlR5IBjNPvfXA2CaeLUH4yNx9pcIpSq2WjPdA+i28DMfuVlQno
cD81uogPBmYp0vguct+UYmKSCIyMlqQLaiyTHce3EritGDznnwEGTWyjwAO33tA66gWpZYXLlxfV
yPRKjcOOwLrVkc/bu2E1cXoLdVEE0cnWCc/kuSys7k0zRsGj3uabrNg+1+zJA7ddTyY9ZP90Toe6
1oF+xLGDy/cPNf5nYwGigGyEUBuCVCOjwPf4gcxCk0dyF28KzJEpt+U2bd/+FoVveKXQvkRzgm+t
7NiFKxi+AxLaUYMovCWb4dO74BmozdHZA8k/EQgddf8nGf4HlATbfjXcfsoPJVp9XSEBLRM7SJG6
xCDvR1sWOVUQkzQYBTh01OqZxWzE070JVTp8eCIPKnYX4LdKeZZxK/20EHbyzSKp8yoc0RiwAs0h
43H36cIxtjPpOF3M8yXNzLEnwBXqPp49hxYeCa40jvBE2XbjO7XZvnueeBr7eF4ZXkfa16N1Cxhl
Yc5iB4LFy4WrzvD3Z9Z7GZcZgXpTpqYj8nqBR5R31R33O3967LBeEsNXgT6onww/4Y8tf1Hk/K4O
CzvlLabi+r3Ju5VS57s0PwwktdY6+zyPcqfkIaWYIalbAsWgqEUpYUhga+XSyHA+h4xSh9cppq0p
JbiLoh237jLFfHSxV5bkQQ1xV8aA0hKnpvjXH7u0dG+BNwrpgT8cgXOHQ9Z1pq23knhcTQyxbiYc
hTxMQ7OsNz4/VdQdYXXWIwlcDnz3wM8sUerdJT0nL2deQ2CXmhWO15EShXkTVm+swpZi+r6I7qas
wACcMJiQfTC2USYGL4Bxpoj2hxGfYoMGG1p05gKbfUXlIOF+8KExwgDCYKkpZbV3EseV1pPS2z7s
dDRGNlxB5nMqnmn3tehWRUeckioPcHoUu+qrHrikalt2ga+mPpdc111QWA2kX1HafT7yGP5FPlYV
a4WhJL6KMZ28/9OSqU7Rti6MxfHU0Cq5hGygmybJqhMaWnaPt5mSZudU3PFrAluOgFcF5X4FzPy+
ItRw4vkRBOkvSpII39EYXH8xdlgIci3l2na85B4WRF7tZu90VxcDRMxw40k8oxt23mc//lW8eBAZ
iwYS7pU3PavN7XIt1zmbap3jHRJ0p9UF70cNJeD4aNtzHkA09V55ymGrvelO/BOPqRDZ6+CwJmJQ
3Gl67cG/oXOo7SsSV0qiqfxsy4nWh1HmIMd6VX4o8hq40IK6RBsvlpYFtgo2YFQjyc76sr1lmRu4
M1JnHhkv0RDO3wQCmiat2YLpTVrbGXYYTH3Jq9XsLyWEZ9YBTvsin/IOkvxZ5wWkNM5DXoN7Be2Y
9CDkrSrkv71AfnV0Sbs6LBvBv5nLuHJ9hzS6JOoLfTRRol86H1BwkZeWkBiTZOcAEYgir44ntWpY
lV8c/wMcE+3HnBQ0s4YwRtHDbU1NOKy6All2wMZJfyfLD9P80V/qtG1yJyGiN7koSIPQB7ATwvaf
p8E5Sc1X2fpoyu17PTGCwV0rZjVDQFHLv4eRv1XC48nHojdLYykIi41jLcVsj8/uEtfS4HvXZ6xf
fNQ4igaAt3X7GHKbF3PoEfIlv+xbywjlmzStc4eIubv8DluaclJMeREsqA+p1PSweOYnPnDjSxug
EiO20gKI8j+w53VhuzZdjkkH4E7L63TfH4tah2AgWpesvuA1O86yCSxL5YL2buPDptcrHVKRcFqE
F3a+pnlBC4GrYQBkqYS6cEeENjunYzhKNLSW0CeRmqyeF4XeOZAbKpvfiFSfqQ/W5yCynlEVefT2
w4CY9LWZLh5MHiPQn45k+o5GHjtETyQ1PP3rrTclWnKviZxzCB1Ewolex6sYkZQYLB/apedy8KQV
IErfLa7w8jeRQujmbsW+SJjAlvLenpvXjTAwWH5yrpsjMTKkk3zekWOFfjONjKcQh4R6qo+ueqaE
YiBgbV1M5Wlu+qPuctdyGLN59/r3JcGqwMLpnKuodsyiIkAmgyL7YRkTLACp+3bof+jpOAhMMYPQ
FgSI2KzeNBAoVNrBTVicV0btdVpyvtWQvmvVBWX8VxRjAafgHfi1ER7euw3l+n+3sCyWioZVTAd2
9s3AHZc+tyAXzvxPYD7O012mDxnP9EwEbqAgqkVDwuR0jhALjaAhGd1DisR6IIYWBcXLEJ2jvwcH
lJLHatJQj77kvIVgE6HAu4JMDhG3eGGd459wSb04aw5vALu+uiv1PX7TeFZ6aMm5O+JZmQgcH29p
0S4dOjGjJTFxEh1CWevgEyXDNiFUEAuInprywPztTdP/QIOqOgyIjkDYzyAqlSdHSfSygc9qm278
Fedf/rUknhiW3fVQ9jI+OfuTw4gKxx4JfFSVAvgwdu7IIL0KUcKD8fIDRSg1QRUBC/KSAOzr2Bmm
X6XEh6tYKagaCfe2hpZdjZoSURmNyWJo0IgadZk6co6YL6bzpQHipLQkOA5D9Uj/YknMfV9c+7X2
JqTiucrw9cphcB2mrTEeizFvF6gI1YnBuP5sl1AiJKt6k2hF7Z0K+7VhsoG+1sa9mCFaF34ZcSWk
oyAumPAvgoX5BEiJqAmjFnF7L3qN5MefTasfTTAnQxMjLfuR4CHnks4eS3qOmwf08WnZG93jaDpw
IOHWuxE8UnfqahTeDR1iO+ktzCdN7ESuK+g0BkdO64PlJvEQAQ3X8dSrJetstLHF1FhKzsbhr1cr
gJRlG7xZ8qkk/D6PBcvYgJXcocH6QMLwTF8111JW/yq7+UPlw321Ee16choaOGYIP87gWmewJMOz
Dk7VYrwOEUqte3ZeecEIgqL9G7wCOA+yQBpbKFsQm05A7g0Jh1Mw4jvHJvob5KETsFaHaax4++8q
ZoySbEoXsdR+q5+YuViaOGf/RRyI2yV6IvfwkmO+WmMXpeObycNEvtNCoWQro4LPOpV355dRyzoZ
dlzKTKyGbwTrKIYdwokyf9I0jKEu+VE8hNU6AkLmDZvfgJ2xoCU+dP2XunZMKUd44J3L8luDq2Gp
D/Eld+0yeW0ga0C2p5lz95c6phzbH5m39qa/LPxWYb1JlrM6tMidTIPoNP+lOMc8cYB+IlwfOMtk
0oQhP/J1MmT0n4T1OWVvk7+sU9sTCjxvDSohuxAehg0kjDYdUPuSmMFa7IW9jF/h63R/0z5Jt4/L
78JdzCA6sknUvQOQAUD+l5a8yesbvjWQZD7bQBJDFxnn72cKB/JERIuSIKsH2XGSgGkauNbw/CXB
Ms8omtb/8Parh00K166gleVK8NT3ZI+5DmVxVW5zNwXYo3Tz80DbdWVaK+rZFq67JpRBRJyITGMf
zfrVx8VJW4kuSDcmpdVYli/4xieyXpFqYyykQfes6SViG851jdmLqFARUzptcmkLwPomKkjAG9WK
OJKij7no6h8EvOQD125fj5x097ORpdHwo4mxRBYY6ge4dINmAsgp0JorMybFu/See6cWJbX9w6qa
fxj4blzcWfVJY0Yu7saYQ2yDHDmWxI6JGk2hrVhist1Jv8lInjhkhGIESX/d1vk6iK2EdXefjlYY
VWhkdNZW5CEUFK+Xl+qcpTeCbz3dAeJ4iN5oIpeu4ZaH2pnMeuoXVmNgjB5RN9/feDwJRWxA59ZY
9wjUgOtU1D0Gn+PBnLKTAuB/UbeIAC5iaF6CP4u/nJzsZM19q96AeZlj1qRlSqaaNX1dz+xN7awz
buz+7t8tQkxV82rJnvZRrbbffX6BJe0nwxAo5Lsf97wv7hSypPLpReCcUdrLNmPyqI0/SB7z9gbl
++g7HsbIBsRBotjN1x7Vqp3gzVsb2QvfczD5ruQKUQAercQMyLTRR3P1uizqqLMycYQ9+QJjP4l1
yAocEicLgOGApLL5vamQeEhHcJv2EU30ZwzHYgG+GKLC9JGQAg4bDWDC1JaFfb+y6P33K2djx5cB
pLMYdNb9CsI5GfUNwcNUBYJew7qXmmac2xCSWGiVKJQFom8sTCEyAnGQ6bOXKFrqvFt+KUKGTBWY
pBxlFM1pM/lYOzeOKq/T/VEcMlkcBsdUoJjbgiCTLfLopIK6gQamQIFLt2ijQHq3C/538xuBd6sn
lJBjIqTxws4OyWsgRI+vipo3kwzoRBlBuCpPMOgjU+y+3+kcLAgkInNdqx24v56k7CAG0kbPQ9tX
GL9L9eHhyJIJuopTgX+1S/S+C/XfMzhoVRR0YyzHnKCwScMlmYeL6Uj5ztoThpFeknm6F4VI9UH7
ohln/ybtx73QuM80CDLSk1YiOtV0lziJ58Hp8+5H6fjZu/1nUtXnCGdMDZhn2Tb1+ORhODngj28x
8QsxyxyX8UZoAFdZnk+/FUlrHZdnZrGwdFL1xBawAQdB5Pvuk5ybGcL1ZQmjjUw6OWdXJNLB1Iuu
IxdCyfkw57x4c+jFKxmRpCDGU+LEMcUZ4l3MsbepvXv97WQ0xZPacF4Em/m7xGbU+SYxxsKr8A2R
fwSv+YHcRD9lRqF7pLsdg4W9DAqlNvIIE22Oj+od6H7txXzoZYx2i2ULPf6gZRjNFwUCmKVODR9r
gjFWU4N6PnkReHrCfZy4X+mdbQBix1uvSxo565YAMnXgviWRtyCjmefyO/jxwbpAZr2H9PPHY8GW
UIkBoy6Owl2LoRlUWfprhaEfAhBRiXb2FN3jyzJsM3t1kND+EyCVW34h+W9YPSpYeVoZ1zdVdhxZ
8HaEgRdCANXZmMw3D1JpcRF2vMmxAnDMTahUutvfbtkvQWZHfERfjBbic/YcDaPnBYklvxVfboXk
YdO6CzfGmBB3HyBW3YcpTOzgznNyXl5w5fbnBh2QAoJmg7pBQpjCZ5xaWEBAEdZo+2AwomQt14zQ
I/bGcmhVKydFWJKfPN1u+7/PRdzH5GJ6UXWw/mZ9VtmnMZMYljFNmkPv8oqH77AcyZc0GPMR8pYF
ubNTRY8F+7bPV2MJcDon1r00+RrMgeFv62smkSdVXjzvsUMj07dUm4p42C05SHj3t5k5r9Co9tFm
BMaQJ1IC77HNmkg7QmB7g8J5G7P8rEbjJf0N9ix85hxhqr+uQlRbt83WtJ4aXu2t7i4eDHQ3FOWX
CkxvJEe9eptNDec1+3HJHyDTPs9IxhS6y0SilJ4BbqjW8bJO+3VL/DyyYoTrHdCnTRvl1Bg/o2NO
9CgTW30+q5Unnp2+l/guk1GEfW1/8xFEBTg7WPWy5u3yKazkdUclKReCpUD2LC7YXX/Rtny88hm+
T2fwf1aI7O3KOY2hMTjd0/9x97wk37ju6WYDT9sIwgnPea919VsAsVat+ioNbhFfUeAmFkRaqUaW
apCtv/x0LFYBO+Sp7u0NSMAkbNwgYaR/kAFGRwQpdNTPn58vgLu9dHW459aL0JV9BUsgaCg7Uzst
WInTLj1zRYIcq8s9nrf//swyuk+g1r5MtFRiHpPbGLDHvGmaow97wGVY4l1/GE0l+RjuKWrdBPec
07K8XE0Iob/TKGKZOEenwedEuJAdfMih4t1yGV/Bz+Uddg/IHY+5cotOCe7KWW0ERte6E4fTXp8d
EcT3lZ0zcfk0Mk5eJP1DFrt730Y3K+72mjroMDY3qzgPbDSQyrgqnzPgOpHbBHf+zokCx31nti6/
zawjcLcl+OOQdrUNRy+K/vGGXT8ml5cgUigdnYNRQjtbpXPvwaDkzyR1qjEiNPtNCyvlG46YLuUj
yOrRgoX/AD7UJ2REo0evK6vuqjB78BdoirCcehUpIvgw6QyTDguiuLJ+K3WRfjfThM6+ni05IpA6
y5u3cDFLvvCVBmUNkjuyGPLVUcswF4FZU27DtWnUtULJm45XUU3bYVyW4Ori21sFOoiQqZWlnSLK
x3irwbVtw1bAROqILcNHuC2JXCrhbEIiO+dNwGOF/H/V64wVkcFKstcTMnlCvL4en6OJxFDeaTVC
GEnSB8yzZvRxqUs8qnDFGOYyYsIrAPZC/YnfTgslUoigHVPz/YhExoRvsuvsHL5BuZHEjNBIqmsa
AO68R/eFaXERyEaEJncG1aCgZupzxooOMJDBL0lTcSWU6jmFXCUccltDTdBYRDoP9GfT0LoeooF7
xgZF+A/Or3y/bx2hISWk0Hk+i83665eaY9Jfqn9uqCJQCUPCkmAasJqyq7Lzv5p0YAPpw58Nwmv9
MOL7qt5BD/l7CEOPINOdF5A0235XUHLkbkrBo4LiZ5nEftzfHSsLrWfg2f0VvnEfXMypwAzYSkJc
+sxQD1O7R79RrGThvgDPh6+KZJLbsmVYs4ogOXy/nqr6FGRzch6HX5r8We03Khl4LuyvydvjtcTL
azXFSLyUZEeYxnec8ILQIaoX6wsehqsyJhDpDbWne4vLdOuM34sG2f7nSCAkJlLSct2ObVuwnK9L
pByzmxGs0cHtwKKJyfkc9e2lBcqppsKv3WpoDua22YkPSFYlIxjMPike0s38Hkw+gjxPRZEipOu4
XPT3AZ8Td0+LYKnG/NSOEA+ZMPuhXlJNywRZ5cPpy8OYDx+LNSmkgTpbNwhglKk8ZBwZ482rc75z
u2Nrt9aJC55G+L4emoAKR6dCXUsS/gQZUah2WYHOXDRVLEDMoo1bgfNmrgdh7aaEHxqK98e2cj6E
SrMnK6SdxvzGohqllIkNQ/ksVZKxYhJD9Ll6UeWULRWXQ6Ibv/6a4EczQsMO2syfsQklzzXiZMQH
YfbTOjr0qBDxQMPlHLDHNXI5Owcxkf6ygMdhzfQ2S4OpvTaHlyYNoqx4OACr1WwFefBtM/D8RQn9
8a8H2oTGRJWzn18EsQXCkdC9pkKJZJqLTyeQD631GCzrnE1MLwmutnaG0VRUWuSRobsKzq8RnuKq
Xw8lM/llu0PqgkbWbLDKGQq2C/+PyVmTi40n0bal3HnEQhCtIpr+42rb6eyKtKHi5BkXgmaXKknt
V1bb11qp7ZbxhL6zG629h0eriOxiwo0jqZv1VyMQ2Gtk651ncjk5ip9DWPwlxFY+xxhFCUmNojMG
W1b+XZj+DidYFYGHZZ/aCgDN28VM9SDucXGFvz1xAFuVAHzDmpfJhN3oAqrp3Y55ERMNBWQoQ0Xa
gQMMicC/jG0K5SWny10YsqQt/MQOATsmAM7qKqqvxe42zSmcVOS2c7W/+AYK4WPPtKeSupmU72CO
j1TUkpCBtbBX3ReJPoQPm+/QVOPUGahRULlVFpDnkXKEowsKLCSrM4LP9+2DYEY3L0R2dfRc0qqr
NJDcmYKJm3Is0nveZzSBxY55aEuPOAEJSQodl5bfMeBQoRWq/jZZJOdHB4o19nE7yL8SpdnfaTVc
8S9YybYul3Aw2YJk4btCVLRpXj/VuWLP5npVSKAuvwSorolYRLVoJf+a4VOdTUehf4nskFTb61Zq
gsO3Q5N70hXInKs67erM2APVHvxiSVzcYRfdr/Z2zqjtYBD3N34SW0K3NO3x/iaKH4OkZCdj70sE
ph3MXhOaK18gIxY+PgaP1OLhKsz2+v4+DpKVCLlrvXs1F/Ysd0+LbYCjy5UUxCVulLAgRO+161Rq
k5xCjFvBwXtQ/kGCKFOz8q91wEKb1hitkyOecqIRGvAb7HXYsr4nAzLQ6XkhRkejytfyIrcLBMoh
Id8huv+G+7MUbisaCtTYcSWbq4Nyri+Ac31jNlnQshQEPe+RRewWSbRtfmVac6YLE/uR6Y/PhvnC
eN6pGzmfH6h4vs3wFs9GSHC1/xSNBgbHo0ckEWUzapqYLFgFxG0gacj86uL0AtC7rWpWacyRssvp
5q+gEYj5xVhXQlY2WBK/UvCNrTgtBmfRMU2QoVxQ5OlnELhcOm+j6wvjrQ8ywgWRI+XXMW0Dhuat
QSlHRFAdYBM9xX00S9NINPmU9DiW02MUNp7wrV0s4EK5aXEFIUrjufFy9IdhduZW/FcP5vQ0Eajl
Ku3P54A58+/c2zUFEengdQrG1oLagdR5D4gsqrmkYeZ8pePt3z7MHT2cqifab2PiHXY8Qjr0rOyQ
MmU3ipQuLyz685hBvknkWNQQbPx4/egZui/wg6FRoFMv4+i1rnN0xmv0AKm5VFpCHkrhaanEwMET
2zmfh0AJU1Ia+0ZTQfzwQdYyqwmYXNbbAa/HU6jGp+545GMLaC8i4qCocbfPC/1zBYFHtQ+GME9B
ltzhjczCruPYzUo7DDkDzxUvgjIydt0fAcOc4pvOFqWQ60r54lPOHTJXjBag9Qb9d0AFKz2hekPx
96Itb7Q52UXivd38qYvbzGjo9zBmSq1UutkMo4coQVeXKoRJOfZt6xk54mZpnfXs86e2/PDAfkaz
r1HX8O8HFLs+BQLO2WvytHmmoHPSw3mc2MRaV9lHhKP/aa3AA+QYoyrHCAZlFMO5R5mkFUN2+bRj
E0w1paP8DLR75RwV3D5IvdcJaJOQ/FFdeUQvR9uT4BTNC1CdJBv4ePcn2PABgbdQWCgjqlT2X7b2
CMn6o3iJpmR7ap3vNINiJL83ZpjWypP626CloxXcOIN/0JQcLHaEweNQC4wlKHjX63EYyoEbNp/y
3v70GkluDLemSbjux3JlnRdYtvSqK5ojpnuNwxtQ3gZ7sZ7FFDEuyDeQY8zcXvRpdC3ZwFXBOcfS
IAatLuEcOd+5eb4xuAplLWdNHNKObn0MAy9ITI509N7c4OMmRv3K1wgm5fghoGj3tJYDBpT9E8IB
1kwJVq02B9JTprBa11QllAYDoa3BIXSHYV+VdrIq1Z2kYp2g2B72D/R0eKsdYNfeBPQDAuvK5Aht
t2VmZrt7B9TleyGOIo+PZvCQtoB4LTDBiJrUAK0dZs7FdKwjPotfRnGQjzR8NixNFLBVKvl4wHDg
NcETkGHh0Hnleqq8Cm6ajld6uqldGcdQzFjCMeJzYMmuFK8CYhBaFZsBDuyVTtQh5D6dIre3pb6h
LhkWXqiwLo2kn+XTmqfXhdSMpnQ+rXiR+gwxJNPZ9MFuooOEIuFF5WV94mMrWIVqbhj/uC/yBsRL
mfyFnlRxA5BAsmRLId+P46dUjdxgv5MEoVXXixQ6jA/8EE0bsJj8RmEILrt/GKiWgc65dvfuVUsT
YI3LptMGEq8SUeLatdyqQ2pTb/O8YMsJL18sKmPYiP1f8t7na3sd5k3h5MGg+isGC20pEedAA/vt
NTYMwhg5J2RgAXfAjjYDb+XPTYCk9hmOsTXpwndb2STvRyFXq7ieb8mOD/u+AaFa53MTyslUzTUq
WOG0rlRVpiJPLALJAmVhqwNlZdjOqNdJDMPJ8YW5uPal3eUHUhrjZhBMx8Zh1WJh0ndyZdwl1pD1
vBdV+g1DEVH6SWJnXur+P/2C1mPV+/nGTnIfYAF2qLvIkx3UztlSVUTPXNiOEVsheGSR7yIFHqoO
ldpQz784TsLs0E9JlTEUvBNg/ccKW9wXRyWB2mRtwxht/pdwiWpUjDDAEoG9ZsIL4kfqzuwQP+DN
jp6HSlrqyehDAgo+LQWJ+gtATdq2fUP9j4C3p8Jg8wtEJ9fg0Vxcv28dIEUSfDktlMzek+bjuYqU
C5qgSggl+dL6XwcUngrZTCzsTOtRwpxAg+VHNY0N+O1YA5xm7bIysP80Fl8SoUrxU4U7ldPzmnoK
LORrSsw2JM8ONeAeSN7IZgQnzN01ooCo7VFGInQKdXTiBvYS3bXWE/xnzTPwfWKSmluhATK+zJVD
MwATcHq2TTV21RZchxksYNGuXwm+G/jyCx+8/Wx8rTLU0ddKFKds/xnT5x4fmDsx+dSbhp/QIJHP
mJ+pfggjFM5bu8VQ0EDTcDGWFJ+5xli0Wliscb+b6EQOdCVZUUUm3pM6zUlK5F4TTTA+BBQFPGoa
ddjxIdNg0lN04GRcNEY+hg/4mOEQvcxpVt50It/wLFanx7xkfjiUSgHiV9ZWFHteZqGmY1nxL5xF
J4cZBBYPLvSQzDnp91ALbQbNPIkxrWxiHEihV/OSB2FPvz4n39z0WrHzPpXFzchmJB8dEo4OPYiY
3ue2v+/XySfhYa13kbVpcg6WoAKrxHvkx5iDbYR4tyZ0SIT7/qIJvbhUJJq92V0SlkayXNS+pqOi
VHEdo7Zzh22ELjOM6Vr19QB5n8SqezBvH5yt71JO9q3YAVCKc6uuaTfe7ArQAtDmMReGQetqeRnS
NlVlEo++k5Qe3hVOtJ0Qu/NeJa63o0EpunO9b1MByVltDkunzuF9iPWy9VchqSNwP7Eyxk1rS6lq
Klb2rQPn3SOfCqF6m/0wlQpHQBNTjBTD/mI1ToohcoFizLHe8mrYR2dAYaPwgUwSiIPukj5fFlFM
pbcQUMVcqRFs/02mnixPr6SeplXUt5WA8M3gJHM1SsBWKH1GKssTKnFvh6ZB/fIQJYN+peBtxpsH
vrmiiNoQInvYXEMDX9Jkf3HLIF4yWHGYw69/DFIyPUBzaPdUy2nonps3XEZZud9v9xR78dJAzasn
7ysvtqiXPjesGYB2WFCD1041zv9aHMlriG+yVEhM9zsv1CNRUIaEEOXTs1HYiXoRaITH7hiay265
DzHTKVH+M4qsDgCiIM/MFPhW2IXMX29rxEqy1Zjeu5gHK1cpsYIli47LKnyYI4TtH6SNItmxXgb2
UlveJY0x4U4844M7JstPcgYelLNRGRC3zP3U15OYB8EwEn7ahr+sVxNjWI3wT2ln/eL0LWFxzbZy
iio+Hjk2plP8jRYumSebVOBTEfU7dyLTzhCfzwpy3hLiv0nPeo1RMSofGfiE2XTLFQJhfSOpLCtz
uoVV9NywnXs/V9brzpQ9Z1JrDYBrVIdQJ7qfiLTmUGB5vMXskYPH99z70vDEBisnqGXy2oepgbTB
G1+QEQrFN40yC1p3nruXzwT5OheUE/Vu2SAt3FQFQwQD5PfGRvfgZc/EFMAnRm44VtifmAQbeAQf
aRghQ12rqZfrljcPDYeU54rxzKtYfkY3Qm0voj7tMQVdvoPpJQ6j75RdFRoWhYwze+1FHljuLnNz
+Za4pilMLMV+lU4shXR68qgOLA5DO4aBGuV85zjWVBFrOV/YIewX2h7ecZ6UO5qbNh3HYabFsgjB
Q/TTMFVeIBc5pb/RiqZ0HDQfnR4H2RRpJgeA9biCP5eFz5n9zPv74mEqAtL58YvexdhMT3gp0TMZ
tFegrgNwuyCeg9vH09OErdKz5KF64yB59fQlN/lD5aP2Sh15cQYvi3SMzBn3cqscdSh1BtQoRtqE
+Em4kDV8YTbNFmbzbnMr933ZdjJrgPVV62+d7qWx+1Of52qGZ/5ubE9QRYTxEMDE7y5t31jbHECI
SZWNHEJNGRAvD2H4aY4k/1IMJLlE16FkCRR202KMu1YU930hxEKWHHSL5xKMHJz6IIsTO02Wx/Jj
ECR9EoN7w4OKH/4wCRGBHlnbgx2JvTe6r10pLyvw3nIKCtsA5g5GOEtv7Yj5Eg7tknwNyWXlRqpy
Gn6bnuGctFKgPjdFv3mbi344qPgZYcsMn3L88Yy9/HaNiZj8o7n6AXaTflzYhKfpIjmX1F56IC5D
c2Y2P/3Vj4qTWQw14z31zcgfOWNQKpKIEwRp+Nz9cmTZDwBdT010fG0Ep+Dn4u7XanpFObChD2X/
YD5idSaalTuJvjB2Et9Eakt9NuDp7dgBX35+GEvTmOssIt0WXfJJgCw/T7YlS+RNyC7EOhk+swx+
CnFf51xU2cZRb1jzEpNSUbsAM1lum7A4DwXOaxHrykUUx8/FAmr/8i7pjK+iW7W+eru5dOWi/Oev
DaG3pZFyhpA1MF39mSLZ8RUiOfvCwwOabBz/izpiIDSkSPpVFBxnZVNdeZaDIbdaOXuB3v47nG1E
fbEGiUjKJz1syXMpNNTEWwFtmClovjJvej5mB5nvxtpV8tx0qFS/MwL+gA1M53h4qTX0cN/F6D07
d/I8M+Y7b+a5RKM+Vv7kX2pHC9aS/XcVEfCJBC/91JrOQ3oKtfQmpSN0VC0woYuBIPp+aag+HZoL
BacI8TPpy5xrzx/ZZWdpmJy4z+RInPvyVFUOVr9gxOf3yZ3Y7OyIfz9YSlUxdgeKbjvaqWHRHgDA
UYaJ29YoWWytzxjbR800p02HmC9uwETzAKtEZC+2qicqmnoh9r4wPPrBXNUOE19BnF1RBZ5KLmOu
0mbQPpJgL0wzwEz4X66/p0k9/UO/Cv7sGGBqN6jAJNaTuLSxVMdJFKW07mPSHTCumYrBYJ8yOilh
dks3kOeSzHQXJnW+dtPXZdPj7LIRrlBqE1K86Z7RifsyK3so3JD+JcYTsuwPYDjUz1AZQvkT381b
feYdC1sfXntaAsiP6Sl8p6/5NZqX5x7q0RbMki/mArKTsrvZlfN9bdrsqzUj97+KUBdnSQW/hHSf
T5T+TSfLyYhOmxjYzh1Xn0ERt8SUA0HTUV2P6EULrkKBfqdj4eJg0F3GYJVBhKfBNV13maEgt8oY
LkriUHfOeZxrWDfEqAXUdsZsFGprxBqYoxpxNz/3RGwMEBpKLadiayBJ04Nh5TNl0u97uz6qrPhg
Ont+gmPpRf+L2UWWxCoQ0fwMoQrwn5otFHvjjRxyGtsS4ovrehcDTmobVu3j/ByhXOznw9NdZk9t
vxkgQb4M2GXp7BYvUeDmscYSqIt7l1EfJvgF5Kod3zXqrImNav6ELvS1EmK9+84sxy9HV8drXUQg
LjFDk4UgwVxUn5ulkbRVixaV4exnigEKOv0hoM1IXaZCVofvMV3HHuJK/kp1CaviVY8GXYZBkFBk
zxyrmHc5ipGf9v56Fv6MBY8koXnv7YxMj5PK9wR8DBIAa+HQXMZNdZrX65YJO6Nf7Vw6npV7Ud/Z
j5i3FJ6H9wLp7iUGa/Ly9I4eUvuKkh8uBHSVi0lTdWmlHkKcFoV0jBMeatgiOQ5+Ng2ZN4XUk67+
b72cpxwT8iw3/m9jmtzsO/CFlFhyHoWxZztyk1vRqfW7UUXAvBBbXLUeH7Ft2vcW6T9Glvntm/mg
xmg6AJXqueXC5W+VDxp5ImwhkjGKK3+egN9DqYoNXiTMmQeRQUZpXyVUR5uk1l3j1J3gZCkeCJq+
1+apqaxSiD8B8LOkypDKd1/EW4GvCyZRCEkTlo4txKG2MuOqGZbBVu/b7jEZK3PqfDgaopF58X3Q
PtxSGnhaGu+gV1XqpDwM/KX155zHfjxdxS1+Co8rjB8FJ6FRVTM+gJeUQW0JfTdk4J3dFKfdN0NO
FWnIxEja/KhMyQ/qLaTFU+b8VV/M1xKz7dnnK/Acxhc24hPTQ0Rk9lPNaBtTjoRnRBReQcC8KxLu
30E4Ta4CliTGJFQHNBui8SDL0rUDEgJQ7keNVRn4KHuoeo1KUy+1mcmFlh+//nA4xSockigK4O74
/mnXyEAcYTmeCLuNk6KXro7dh5NdXdM2Nf62Gt68TDWX/LV74rh4cwGCSjrMmGW5FhcyPHs2n9Dt
+UfL5gJDLAZHOrTPe5kLhg55ZrIw7nuqEP2j7ChGoPPslWfu7ROCI5GXOuVeu+lF1ZZLq+7dvU7F
npsz9dDLlchgWsbKdf7nz3096Z39wtvRFYTEe3NUzwAIX/YtPMg7UV2A3bJd3ZHTahztCUiPBs8i
StDrkZ4v/FEFm+P5CtmYidFhBjj8Sx2C1f3Y7T9ecny3y5GFe7NH39jiNsP0x2QnHO6TsK1Jq8Q6
iqbHlcXOvu/LEQWpMDr+/fme7Re68TTGewfdqpP/e/AXWnguzOje5JNmNPh4/gr9gFxXhImTcXgX
rrWg/gLeI/MZi1urdbisWXaaJZ82n32tKWPNg/GrYsOedKwx6USatnsmMCxJ+Vz6Akuj8+f2K8If
me44cM7CMyIsyRc2kgtjWkZSaRt8l+08QOszfMbqv8jkzMQPu68169OrN3Ds+pR/NfoOYb9E2Jf2
Tmfr8XqOH2vGxsG40SXyzYjXwQ78AkvF2JLFVcxv8hGyedtvVhgyfKGO0qyGkvv25Qj4jE6xUS5M
/PXUOqrWivYFwpfpjKDoe5g/AXXzluegl7IaSRqiNS1/RF558pyTbndgR9wq1+cYan02eEIDC1Dd
U87kh6smkn5vO2BGjI7v6WlOv5Tr7tDa0Zi6J4fRyQYeE/lspRYuXC8DbwBK+tMXLhb2ZMQOSwM9
a/yQ8smXw/4QkRac0ZjFHmoE1UEp45IcTm5zPmmSSB9s9AL4SLiIyDdih+dmoTxoF/PhqIbx08Uv
5J4ToOv7URYyY4SFhiYaw9pr3zpHj52fOd2u76hpj1FZpuykaKjh01T+yjo3zNQ/v4mtexV2WP5/
dU4hEsV+ltD4j4VL6BZIt3AQTbceEQJAKKEWTtX1YfBG8imgD7/oWZGDwdD20+vT4qIeur3kNLvX
B/19OU5q/a7o54nvdEM1yz8OMJAEwNujrak73+cErx+XLkwqb4heqR0n8PG3wRKr39/GwjHLlByh
D7g69Pb4qa1/FPKOJ5UdRfekiXH72bGkKJqiMQLS2gDLBvUE0BZFvNyljcuKFJjB53iCkmTls0qE
2tFGlS5lK6FkBt3lLGaRn8/xoAS7oKRg/USZY7hc5gScXIG44IGDud50CVLLqC39++WeD9kquBCz
l0jO7gV3WNpBpAq/q6v8FhEq4HWnSlc+jtGgQurZUcr0dQIvaTe2Qby1rm9dKDhqUQzluKzCIzO7
B5Hm/mFBln/rl4gmMGXxz+ahOs8gucDMhrSSO3RQLuFuz3pRh0PQojQe99YnjPZ7oNHz2bdytDkT
NZZSUC6i1tHyBIm61sWghxnlW/zl51D5v5B6zv0D7a9xtetF2wl29eQQ7G5FfGQVvz1cVPC2FqzS
SZXhm+u4NYGTFE4f1ERJssLM+SiAV19EeF0rGS9aQOMx44GYn4E/apWXWTaB29PUt2iw+kWmKa0y
+1JJGuGMgECAuGSiE+4LaLD/RGcLLfLbh64rppxjYN49whniT5S5tjTwzQGAHNW0GOxZaQNC0SIv
H2MsCAKGGUzQmEV6HRxAPrC4pr1nTw7LPqzr6rfCGA7ywrCiYRNfflnMH5md2yiF5GlMviaBiclt
sbo6msFb43/bohxiIYXFGnpPghcUEGdV9fVKQTHfIGGnWXOuoFUuxNGHxeF9OjrYMA21XdkUp+ms
O1GSdCIKC5Rb8zkDwt1lkNCmJUiTZ3JoapZMa+MJ2I3nSvKsW4+e1oTw3GqOTMeExPj4n1bKyvX/
B98prPUsx7n4LfPygBVZb1xPwbAzKV7fQYcHSe2W69L0t/wCQ57zKJDUTAb9RLQuIVjMuk+Z5FnG
wHeWxt7QX3Cup77CFEJN8azAVlIHCUc2HYK8e5H5e/c2N3doCZqHt69zNKccYJHKOEnIn9/iOjRC
AIuD0FJxsYHXyBRymnm5YcgolucQ7rTYHl3Y84otrpOC4cEFttWn+/BOMY9+PMEn2vwdt3Dcac5v
3PWFxTrKdn0aZeaHF1tILUH6W2ghOOOxlrX+esb1YdX+PmcmlgqY+I4A3GvVZCSE02GDgq9EKU/y
J8jldiV56zdtFcNlc99yH01aPX2TQnp0ESWDXhUWL7Am7DIkx3u1VIwW9JSJZCCBsVDliQ+r3msf
WayVux7fSzq+lExlFMgXj65xaRnTzWY62ETsQFK+uHjovx7c7THK8YIStTc2y7ckXgeNav2am4OA
uwLKS+nZEthlVdyeGffFqhZKOTgznb2J6xOy+gTdAdCn9RJQaPW5Oy5x4/8s6eboZIbevt2F3WYg
4EpvYo4QjYsTlb6/VFVxRUvcb/k7dVQ0TRmOnG7UJErp4Hv97dLBA3OEf4sSlG1MHiAtRLqrQz/F
WzEjriAoTFgn9ufJBsIiCtC80r0jwDqe+G9zZP864JvyzE999OYGbi6efhpYQOa67V11yETT+3IB
HQepuHQMEBDzpytrToEoRvdjv6fhIL0dXKMFqWIPEnropLuXwRfO4xkk+xB1iEOU8RLZZTIv324o
XzqORsUJbVoJPwLTrLbQaonTDr+s90i/BG6i0y7UZSb9gC0Lsa+PO4WD9UnuTbtiPDHJnnCOLlV0
GL2CP/mVgEv9/eGh0wU/G3OdvWiYEvGGSyYegQFtrZIexe+nlFQ2N4zJJkYrfW+bkcetxQnRdcPj
u25hh72HK0EAhmhYLdrfRsnKuyjuZvpo4iZ1FH6vR0d6tLznBifexYEuLaPc/kRJxy+HY/YwFQim
sEMcDQOS1hdez9hTZB62AhYxM+kROv5lCrThNgNqEkb71QCAW1d/VUVPjidJv9Ol+Ak70ODQ2vSp
U0f/FOxne+ZjuwkR8Jf1nLQydCwk+4/rvGcOTSaBCRTXEZhHOFHAZIMLINGuaM5oLTOAWJpbSj+q
T9gIwiHPzOEnmD8bbMYGRAA3B4R/+Ec5fpf4cPJbszLuE+Ysfhk1+tUZSUQ3UAwHySMAO2+bw9dT
1IIGdL6uXowbOKi9etPIYRW6UgDlgqwWzUa6unaNiJsM7iyimtRmZMZ9Ld19BwE+OYEL89wvlMck
08C1fw1YAObICe5KmpVhhTnlA+z6Bimq5KNVrirKuki/ebNquyhpCCpEmwIhzFNAOP8ZGlqEQ7+8
jlwyeTuP+nSTXfXAPrehVfrupKHnNXG8SdFS9ZBZnNVNYVnFtDrRtNobstPhIujhktDXDvuYYiJe
NYmyBDKwoL6B3LFn4Nyns/jvkB0R9tIVVQOmGkU27s4fHBRNtPMWJ0iDGnVN4sVNkcFqLLKfTlcQ
Sjqs5WC3GTxSVzArbifNZCyMKAqL3j0RjmKjpJtnw510Apsf7kkS4ZfSZ/R90ku0k+/AYsLhpL3Q
LGQ8p+VWjkpyCt1OslSPllbMQrEwTsu5esGQdUgCVIRPzYyE6j5zTOtewo/fg5/wWSLt/kIItojz
OWz7/9CEdFaBlQrKV3c9UU/YUFUntEcUs1/8bzoKGxKiqRASprsvbYDcuGdt8tTpJzHfBZkZvmZC
XaujDP2Syf9wD5uQ9hpXue3QrV0iyssaLK0CSZ0G648aWZuH0LVNx1NBAXIlzHLQFKv11YgzMzGb
VJc+6q0w7E+gK2IY0wgftIuLmYt9efM0z5jnFkwhN0vW5tjIv6fxcexrg38cDkQXqxUvIZq/ZrXH
jcIiKXmnrioZw0MjaG/MHI+7EXKmi58habz7Gf5ELSkKc0yqI5NHLi0MAs5EXD6S6JlvDh6RRRPU
A+aCehtkLGLFNGiUkp6MAaPPg1DOiurUl8hYE5VwlQ/198XqWlYIfSCVFOlWExIDAgbmyrKwU7zu
W85L8hDGfvZpvNop6NxAmT+iBR1RN6xl6dXf1ekBmZm4NztTk5DvjG1vGHMSXTPfDKrozKnWdz6P
YT7BAJCF2o0nlrVEerWDS9swXuvgIB7091sgwwVzzHMrNEnV83Umkm+sblDdDb0I9yoWybvT8op0
q2SxSx8ac1WepAnOJHOsPrRbm/YlSPPrsYeFiS68tRzw0FowMLFyfjoyg1la7LWOKoHfL2oMrfqn
+qvQEW/byin+VGBQw4XGpXrz/uByFHEIR2QxQwqQuO5QvUlJ7g+TR02eQnTl8HHulMdp9LxWAycp
MxAH5OnF10/XU+7YDGEg5+DkPnnjjfAD9UFcn1sa1euOFGgpw70OM/3ohNy4rFUL3uyc0h1AAPEo
zEyB4/3SrE6RuuK6mla0/NZ7oY2TrC6VxmFJSFMx3HiyMjPrgit+1QfZ0qZlFsTqobf5Ee8gH4EV
paPrxsyZ8xLsMSdetPcfD5uG00FUsWKeal7y+5DR9wcd8Gic1MY21f9ZMzgfY31k/6FSMiAqP7jl
3Axw5eeOrm438fSBVwg8sQhAIzEl+N2O2c4wr2BPEd+bSE7gHhGH/qZH3IoQg02Po4MeZwShlPMd
EMlji6o0jPsiQsXDsYCCFrEjKbyNt2u5G8DRnG4I14JylBKfGDQVLkH8m+w8GwzH5uHtOEQe3dtj
CuaZviiGgitl5KHpU3kYg1PyVjkNopjMz/ZtDyxfhZQgT+FXJydeEhwzaVYgeyzEEuTAB7M7ob5H
7gZ2FjwBFFX3e3+iRkhR5+GN0kmhZi6XRHyy3q8jU2XamdTwGxeeWIRyB3jx1Vxnom4yu/702fTT
2gG+eF88cFFL5q7tMLE0N3TPSGvIB8SeSl38Fd/MBwqSbf9gjMUnGkS0A6NlozN/uEG8Rd9+c7er
qEGDMOTenoihxjqwTlgbZfvZQojf2xI2xhP0d5UGfpCNawmOwZZv/hcHK/Ka5d/kott7TTBVO29c
P8WaGDDntI6YWwUMRSe+joA3Khfqz1Zvvso1oxBB3WrDJNgIdpkIDHmX0jNDzMCUZBJQMROI8RWU
lTQaRloUH+zelxIBEIT/rdGo0xNOjF5SvbNzjb94hrkbGRirr9c1QxEFrBUQPqEti13ckXzFJzyH
/AotI4Jo36hi2s0TdH7VV//nk9/f7FfgZKGf0pp65fN5b9ddlkEwFZan2t/JGwGfGyKUXe3MVuo/
lS7PbTr8g4RM8Uk5ActVTHdPj7lKoEjc82EFPT+puezFEm3fT2Hop/u3JHHDjZiAh6jyQn4t2M2i
JZDqB8XW/gsmHjZJnJaQt/HBJwDtDWmDh1TuqHjWj3hs0kT1maPyRqcR7VDjMx5UZrPYJNL9I6Wm
smytSQnmx4iwsl9Nn1BZqtnZxoUSLEuIcxT8lH6RPyy4t/HoclITiGkkKkKhDx4CQjWuoGk/9A92
yDH2Hx3a2TgnOGa7cfleP2wjftj7vECx6UOsYXIvUysVXhe7vSvLMeicMGzgFa+vv7kZuSEvbAin
OgvzF5tYeDKUQQ4VexHKx2UBfJU/0YRoB3N1Q5OrdCqqr6Tfj8IDa7Fr9H1fDN3vrZ07pVo/0ZUx
5735sVaaKaNOMf5xfCv5R3NlT6bWzlD1pNz98x1/6r9r9GtbNdowPEK8qHKHZv0me3k6N4l3QhhF
h0CIwb96ENWfcMN8kJECPj7WYgbSoPtaBVI39p+q3WEcNZ+jONhW9qyD0FZcoe4398YTxYgO+EL9
r3LzhcJhyytcxr2zN4IrZXwE639CeTmoirk4SguD7jyPZuDsgoqL5ow3L6/FTYbGe+/gxYnt3SCV
V5MRnTZ97sk9Glyw3mvExGbqWAM36ISZb+UGVJHrIL/yVZoWr/gIguUb+tCg1x037SjyMv/oOCUT
86/dCj6HOYS8HfXbCvlbg76bMZsFnU6TkcezAdRBnmyabYGJQJKP9I6SZfOm7Wd2dZ0TsVaX1u/b
5wDlmxibFqW745AhR7ipPSkfyYUPdbuHe0XYYbMC3ji7jei2YmhW2YW9yKPNtPq2cUT0UoN18wex
ptVX6+Nw46agcQjckXTd/ORkJTjJoC46Al/8BKiF0F20CFSc7n9IkiFqDCpeN+J50x5BR+OclNED
CMa+U1Gf+mlw+8YI6RaGQuEycbAnBy/iajPtglhU9FblkwgLClxwfrIdahrh2rFW737XfgMKk4Au
3Qm+n3TmsGp6h3mLEqYixYHmNNJNA/fQKFnhL0kgPul1YZSGETUuQGuRA8oH1uuM95KxWTWnqcAT
B+8oIBL4fqXiQptkxK6vvVnYhUzouTeO/0vguWZeGWe8sIewgzAoC7BxbOj2vbRwmhMI85XYKagw
AZOueu9wniqvsLI8hvW63YP12IcAkPSQlgVovXjEYJfBwNqAEFqAzT1QVxbQz+35RvRUbCj0YgOW
D0UFH8L/s9/11ge64RtKTZHn4FwsyDyQXy2b5W1HYOq9zRuZcML83kMQqC+kdGYj7H4sUAgiUqT9
XItItoTJ8CrbfSeElFwtAHW/zBs6ofAbyk3bDbEXUj3k5yEmRHz0K/VFNrhM/ZNo+Jq1BY492Tv6
hUXPNWxduU51XLtKU4k2fCKt3FYVjRbndHd/czN3hnhcHnARZNy23m60lVdBG/tuZvXT1FtD2UBi
S7DMzCuMkgUukZa/Qebg7wjjWxe2vGqJvBxsFXQMhJHezDTlBuSbXdGqsvf0FrPaoJcG0gpl6leC
Nh2qlQnDAinjwtiYOO+AbwphgXSGAoXM2IE0z5bDRf6RVc+0dROTs55r8HVhi+7Gtbd/vF4AT/B5
X1S8r0QVYiGVFKO9UtWP/S9yfe+hJtL4D48i4W4lYvx+vydSQZSvygwk0onHLUpoiDYQgeSLWR1O
tvLfgfXUbwz+jhvzhakptBQJjmCuS1Qh2VCHlZd1FtV2H93XIsWAiiVTpV+8LvuOKhprb+Kl5SM5
UpnmXuP7Zb+1OVSrYvmQ9pt9SuGU+1ReWwM1tFSpsSETeFeZCupm7U9spmBdwmDOLt/iLdck2L7y
pqL8weYb0i6yQpz4vp+NeHIbpLlgiYp2itoIBSLh6K6VwjejNDT7nbj8TLTtK4kFq8vz+ljQ1H31
Cfotnyb9XI+W9FumKAnuC+ydu6UMj0oYTE3qNa5t1G10jTpfKVjxUHKslYzEXncYRleLCNGisdQL
Z1v+oUiZJEsAmNTXO4jiCuIUCwQqX7DEpKCRviM1oH0PMRXMDj6ZZBPpHtuNQqwgBK4IIMq4QfC/
7DKQR7UQZLssrCr7BRMtEfwlEs1wDSk+Dv1yFMASNk34PfdBhGk/iwjmpi9og3W2UmpztDupOsKV
SKNkft3xnvzBfBvOJWOHaN3NsMuWY/0U+KwDvELl4iRDTaSKFkCMTWV1HM5bjJsu+lAYM4uh9EgW
OAb8p/KlckoZ6UAR46AkmFLk3LcHYXupQvsVbFI0Lub9a7aFzkTV78QnNjmEdBzijmAe9Q3He8Ry
Y1twTKegSbYknPEj13U4Y4xSfaCNWbB041FiTvRmwTmjOcv7XnaDQd2/FEQHFufGjif+oTSyV8oU
C27XmEgLiiu4rbF7BUtczt1C9X1fzhoUMKOql9VTPQalKSgxeQKFc6SClXhUdUtG0lLp08daAOTo
PXvMSX+ULhVoCFZG3I957g99WypsLOBvZZApQWoOfe4Mke/r/KxRmtwiJ49OKwhE8SNQth6COgU8
eDMUF5I0nO/+rSatrx4MVW+zG3WLEw5VX69md9MXWsPYUGwhS9RoYqcDLo6u7oUYbVRdxnZTwcZw
H4qg4akksC//HuC3VumleARxVIuYw9lr87n3R7YuyXhIE9RoUtRpsf9LELuJgcJf+iBonFcbxc+A
4mOgoOXx/ce/z8kwFo7RuAmkAvGpuQM9GtBvV2pt7EqLzn68HX9uvmrYQoee/HHCfDMj1j7KY7Kq
PMmBTRCDQGV1s6k/y4eWGSNvDFxQbgrEEvrt76MXBp6juhJ5C3hPSUP/BL1qgeMEZaVJ0R/tzGlP
LAvOp/ogCdjUMnvEAT/tt+7YoE+3H70ZSlqiYGYYpoJsiDLUeWsnGyc6lEoGLyX4cZa7zVv6v7bh
bAFzhXVrow1IaaWgd2UdTXvj+oIKcffyh2PLc/d/SGGvilKatJmVqXVhDni5/IQ+OtrSyMtJxhJg
5nuqHOodV4AUjpeqbUsL5hNrP2uAQA9IASScr7KRQ3yioccg/co9V3CwXGKkjMtacddRZnoOY17o
7ZuBWT9HhPH9gjItwjwgM5ZsWbLiv4PeDgIoE1Dv6V7c3ycTuwU8UwUuWFbR05PyluVvlVdL2hHZ
kQLPo78B5KJkvW39njb++knxhjWBY6Up1JlycVazbN9VBq9kbwUfQNMga9xEfSX8u+xBqvycFcHm
y0QwOk9jyXB0Rc71BWmmy01qoT6BgbTSoJPbYcyFThfIeUp5GUzHAWfjbzt5f1P3Mp8QCxgk/NXW
3d/cUT3jrtO15so86S2zA+pvNUqkDIbHMCoKMsvBwYPofFSHnQ5eubW6htLG7CkFEWoOreyHscUp
9xtL5tlwoP/FhelwPMSphEzKW38qo4OU77LbN2ibNGUv/MqXc8rCPdk+n34wI+TkIrTncssgQjTn
FVWq6ayhaLgwiNROFqKMkHrjOS7JqCUXr7OdIYPfJh2Vg1t0+eXmFxqFa5lo9M6meqhux+PtE6pv
2gJ6AaoGQwgq3pvW2mKTv7EGzOjfOfbOUpEIEhTHT12d5wldXXEtBvp4QnfNl6HZGCWFHQz6KEDG
udM/KOo00m9WnLR05parv4X2r0WEUCgBXR0cdfM7GuW9fVUnA34nc2q0hM0HYM/fecfpOo5k66/b
cXPbIKXrqbknNQq40goTnPZMAEylpckscrq4PRU4AQE6bfWzf4AmzXxon6PUuyQIHMhq9JWK/Y0B
fXiBqz1GjRKN0uf1NzTpvGW8GwmAL51EavjHFpIB6gC9OR/kVs2Eh6+9zjJ42k4+yEkrw7hUeDUq
/HCyZYOJL7HWUsReBp+4jDb8xOXqd8q/8DH/qtlSYQ1iz+6fMlntnCKjGG3jTbxVT60Dmn2n4P3T
b4dBH8L9kTAjQ1H/E6VqGT1bUiZrcpKdZy6/WdzxS/D8duyfLVqHFsXpO5I++Uz1pcybRhxPg5pH
ItNg/EFW46PmWRKcJhj56QXcE4ZuMo4e9v/o7ESgMtiK6YQDfhMCyyBPrKSVBi8yj1Pj4TnXtj3I
AZdHUYwQVR4fKNLh64ZSMOZIy/y4UtE1mFPm5pyFYD9Mz7iUwB5WMClrZhCtGAtrEyJ71vWra26U
+YPp5wKa/BzbH+k1rQUP9n0zVpxooa+a/oxS+UbL9NmwZPFtgAMD93MJTKvhbAwlPRsWIDwMCc9x
6qeDzHCCFJ9mSmrbASgKD9Extut/KAIDP3TNvw6dlH45g1ysFWNStgG80Idv7REXIb/GQga4S3Rd
O54PX/bq97y5RrpdOfx58XW4p1LgQiO88zYyTUtBp6KhYdxPEwoL1sJ6xgwlQA1Pl89B0zgRoiis
ad9Kp4PfzBCZyKzciYASY2/lxexAp21eimPyuJxsHb92ffz+mqKkHPE6xAto9jvMoSzho1Tna5Ks
AxE53iF1g4uLM7W5eMNHQ3RdR+J4Let4h5ML6SSNLM5MkRKSQ8cPSOVLGT73/X3DBkSBvgnlMz4j
Dn1JD76/UCbcuIsSTUeJWWnn09OqTnvj74y5ksB4ccoRD/dx3eyWVRagf1VVb4PgzmpUfWgzfZgu
mKvBs+jew9oZ7mBf8tpPuUXR5aVNBSny3lAyprkHHf+d894DOXt3e3MTfUz1dapiSeYv2S4f0q9n
6ulWSMniuHKNvYFHBPC02Um1a5CZRyX0noCQnFO2p+MS8dcFN/XflOjDwQ8UmJ494nWVIkAYx6N7
EJKTNmkLNsYpaXKDHaVMyOXB+6nh8gJmF2LzvSKZjBEiVi6aJZFQ9mLoiadnoiAIBd2BcAByRj3i
8G6R3aHdDZQSMkSxoxJZL0WhDMYMtAYGILoge3nU45m1j64d5zMjszNBkEsJ0YuzvP+RwfA72+Yn
MWbdUSOyGilcZ/NRlE71Iu4DnGyBy1h2fR8nXemx5Qju9AHvaaTtItYucYWFSB6DEDQA6vscWhnw
+y+68jXg+GyNIqTWm3NbSX6viIqIhoNYoB4ah0vAzrZE8SZ/xY8myH7StwCKhLI05o7DQ9ZqsNx+
BThbm6LadMRZ1eropMq7KWUG+1+liY118dofKi8S3k7RcSTMQ81eABGMdDsR2AhYpn0uuHtR7qqG
EHWBjjIBKnbjXjO5G50L3ZwLUwyiOglLhwsPXXBTs5Ct2Kihk8f7IYlmhudyrjsnXbn0zYgPpoyJ
RPx1MGU77QvSVfG/9/6OROFUtrv/py8aB9mY7PkylBFakzXoolxtatjqOkhV1EBmuNckkmMEp/73
VwMsL2n90XDbWIlmxn56ccecrZlkQVzZPAE52yHkcChCK9YEGTI4wI+TzpDKWV74/s1onZat1wuB
vuAAMymSbzuzeQVk11a0qVLEd2haWQQaZAZWzgSdABdImBwx9ZiSpcv4c8crXIHDCZxjfCk+Kg15
iIvOJ76sT++GzRR43eI+6DjRmtceokBtlXkJQ/F/Tq1/oRD8CXTK5LNHmWJBv9b+LHpXqveeedIi
sPyU3vJxO5Wv8ImTmYy3YSHB/p3pq7VkRtfbwn7Itl1mPCHLAjR15enBseTvnSW6REyVo/Sc65id
wHq/eMuhIAKFxiF3YGFb7m240w6DUyJosyNwIVjZ/VT0IwgLz9QH9ekxHAeg5onh0w8owqhFFG06
NxGYO1KDVDu21QvlDQYkHXSegnFnhMoIxMfF3MXhXwatEVBWUwcyUJLNazm24ChCru/Qv341PvwD
Z4KReGn+YUosk0Ip7fjwXhZKTM5SIQoyjVo7QfxEfOEjl9z9yfYnpbqPgCNQKx50aOyG58BkuacS
jwcZ2XQSAwWLnUYvhG6OdeW+4xoWu4SyT6N5RJAP+SyjtRWL2s8sWATAm6scLbq5XqpBqhvbI5tX
itC9Rmo1EvmB24rCSRojM0nyFoqaM+mjdtgxmZO4s7iSjuRLNt3mhmyFt3nD88i1YCoWHk61lCiN
s2sqvknBHiPgq2Qm136HJGkUsXMs8obn6nvXu2EjJgwIdX0gHtZ0M063cb8PTOdkO2VAWYOGqjXd
ItYctgFewavIzjqjdhWXC/d1MHR2tlUY3jfdvd25KxMoRxCNy8SwxETVcR7uCjKBelFtSYYUX4xP
H24WMA0nSbzNlTI9M5PI0cwKGpzs60kGCT2OOgv59HlmsQSsmZKnhqICSSSCD8P+NOse50PMyxMS
bLmITELs4gCHVplkv6dyaZYMSVTY65h1S3mn0d1CsDv5id1tJBcHVnTvnA4KuLRnCu61SvtV9j6o
AT4IXTKEJuXfXeFBfqtUycU2RrbOaFbJYJCSIoxA7M+X57KOPNDdbBDU9T1AxPZqbKnLuEDH5tIG
J9g2TNLmQwLpV12dLcPPVcYxUPjp+ZJ+ghK9gF4hsdodKuBzX2L/CW8h2fwQoUp1rJWnWslW/GdC
CS+eRLAV8i4SkijxF3V00WoTCYVq65MG3tHqV8juiqzj23aKm4PCTcX+F0WhckUXkf6B/U7E1W0R
2K2fnirQWfriByTfga5sSkFcvgwOoHKh8ZPAeOujYMSvApfEx1hp5QJmTf2pHHIqw6R+WdE8J0aV
c1sLy/JuHTiHkSAM6MyktWjdDhCIZMsHE4M0zYZy3/VlvU/slFuklBmTpS4fjRMS0Eq3t+81Vyke
Nz0AClEo+6EQ5dO0EN8XNhSRnS48Xv6s+/nk1L8/X2hUFVU8tnZe1BhCQYToZh0DsAKrmvOQDwBm
ugeIs8LYNZqkT5vgKJpPObP0mssIlMiy6CJik7cC6Pxjwn0d7L/W4TVh57FH3s1MMheZXY4r4JeE
jTANjTX2lQcDaKyplChuQH85NLz3vECbt/dIX6C94yCo+x6aoelg+Q4lwmSakLz427mtN/J7My74
nwHui+OviyzKH27OtffJUMzP67g6X5IFlAM7USPuSMOb4h3DxG2RZo+q0CchT/WaYBR+6EZbRHA/
xe6ahMNrNgiEq3S2kDPoQfbpN80azcck39bloJRMD8WlN476kmJ2zVudyz5Ydjd7bzmUQuqEIWjY
puLkSj39AOptn2Sq5+ms3bxY5xJ8DKMmppc/iPmyhS4FzVzQ6dzTXHUybQGngU94DilDs5Y2JQJc
uxPLlR+z5QFbQUA4+PNBkmxlsHAiMtByxMkygMH7UvaHMBrToNRa4rO6vkecJ60Xi9mD625Di2PU
ZX6/FHWSugdSXhMUPcyGODV5nFayiHm+WL2wfEWWkx5riKhvOQDsX7s4CAFiUeo5REPnlu/+jUMo
hXBiQAP9xKeqVz/zIJcnZjRPZim9akMPV4p+8/w+uhy/Uu4tN3qyFTig8+uTu7ITJCSJ1TcV4kB/
tvpU6Olrc3+LIlcZ+EzyMgFkU+3t5WDs2Y/r06QLt0b/VxTQhbrI0KDinwkReE0+hhyvLZcjk7LS
qlw02Ow3Z0b1vBUgde4YVf19nRyF8FoPqiL6+xrDxzETuHrB3Lg17lVlkcW2uZsCnrMboNopaGxM
C3E7TqW+sloH1MqBI7sbrNm/UzDuTfpS4JGFjgKjEHUo3EpvdjZ3Vh4ssYs7qlfojcYgzmHampka
RJA4TDRqrDDZEHFbXVbI7ufPDAUGd6Oen3RvAW1vPLMc7SVqkIDruBXmwafo4881xUT8wpwhrFCa
pTNYwyaC+tZ1SZ8NC9WK8HBMWVjoGK6tE5wxZOdYAfM47z4J2VzAE0fWF2umsL4M0fpCbayyn4rU
1AsopWBIuW7HZhac7cnHsAYJMrkJ2sSsJEw3hf4w5E6d1aD8Oip7NNoY/Ql1Q1v16gUmFIw9vYVX
ViXT3a3u6O+LcBhxLAgm3FAeeWDu+t4p6jtbLLNT8hOg6H2EpyvRg5RFzo57xlZ2YOLY1+gjvOWT
/iv+OfXhP9DcI+QNRV5NkUD9Qacwfp8YZaWYcN+KYT+vz3BcY6bgi/KbdrXB0ep0ihhVCyZQ+buD
k/YWyfLf6nCTDMaOyASVscecm1qm6uUuBe0Up3eZmaItetfHhcCQjaxFy7CV8mQYdzW127zFpgH9
5SYX2i/igOcdHZA1qYkLT8d+cYYsdB9C1OF4liuWZDFZRjZ95O8aoDluifgbbPuUNSimy/xsLMhO
43J4/fwpmtj6AVpigvzOYsL0zzh7XPzMUw8UoDTtkJMuFOfwJ+CcA9YbPi4iKoFCZCxhzQTwX9Ct
ojJBgIyeJ6aVhtb33hFJMb1W7evU6yJ0fe+KCp6pN3aBvntTOQQlo4E83rEchmlOhNV5PvNFHUSv
Q7eEh0EaypgSjmFFj9aQKuWNCr6lP2L3ObxNjhE5Wo2+Gug5a6KxztN9E92NJr3aBu/yKPTBmVOK
O8+jvD9mz696iHEvd/dlE4qqvGWqltZOU+KpXYnJDWQX7nkTub02h5gyWuI1igRvSnlt0hskqMuQ
c8usAF+AtHonh4Qo4zoaT3mbKZaiszJfxwGUK+px6ZDNtrFi/XPMA6eaDPbXYUOmGWPVbOs8rWTy
0Sjlbc7ExsyicZk5OxNTGn/wJ1kyHtg2AqfaHXZeVyxC/r5g8rjZNiTjBMlBYzXhG2kMvxFN5sMF
Otf1875d0RDhUwXP4z2s5FvArPtP7bW1nagNDQ+Pqm7lFk0/st1ekDrDZc9U4dPiHYiex0oHtCf1
0NOfE8d2RqOcmh/puSwHdPSZZfHSfyhNrpWbLr9VsmBjfC+VRAIFOQOxUrLkgOnDkoyNrHNKWeFR
g/spVLnXAp0npw6UfjvXO6vhecPpj6r7tpi9HyHG3BXabSfVZ3DWAax6DhG17MmYX0u4Zkc5Aetc
XJJN5dBn7ybZEaN1xDmgLbT7kqukBZgKC9R3k5qTiOl+NRyiqerOaGLGCYag9KkYh98+41l13zNd
aeY2D7u22sf81LuslPKA8qUu3YckhyeMXMyX0BY65NHX7OLQBXYmGgESOcLWlvdb/xj8Hs1zuZZN
VLoUkmBjn8xNjuDB31Cse7ZBuS55SX8Jr/Y+5O21MMTZmI3v/ixHXcznW8pCsNeOaMn6P6m35gCM
TMJaQdEe+Uvj04VL7n2F/w+qGOCIJYJ3xzNNyWgtNUJlxxjAGC6vFIaSYXyOIuHx+4czwQzhLwQp
1pq5YX23hjRTolbKm6E/myDKV4LirRDPXfTJNO85Mf1OOM4MMcwupIFAngX1pYUJx+F4WVJYayqb
OCqt82vsHvW8nQAjx31JW7gJ40KhBg+8mWxWznPMqE0CYi1xL/0E8gK/cgo1NrK0e+bunDFdx9Dw
HU9K4zITdc8wu8ci1LZItf02du2NkO/GrYYQO2Du4U8+ZzG1B3k4iJob98RnYNvwjpfvjC5r6+RA
Tzyl98to10M65pWZLRNStd1Ydc3VXmzq7W76dD1ssTCjnHEZieBwirg9qfz1Isgt3CnTN1Uac6b+
IyNXElPVwLguiO81jYGCGBuVBdkugdaxkBMLi0bw6Eb4bV+N0jvQJuLZ56urYP6zbTW43UCocqvq
7NZr9zG8+PGxNvcgBLjswNKBagVyBpEdu8tfo5iBSfHbkR0Kn5jz5kdw6CThFZPk8LYnWUN0Q4Ly
GW5GkAXaEPxCvF20oAfqKe5VDfIMyo2dbbRrNFWrxMLVKAFqiVqv/+qPww2ESNAvitq19hT4mfuB
d+amgzuJTAELhEgSZ97lljywBMlDBtLjHMlMjTf/Up9ZbImx6XhncAF7waBantRV2QynR/io+xtd
wu6yPCTYBg7weTKsjOOgYbyyEIoK4ai6iwa0NNa0+d8SvSJzm5gcS0Hv66YP/kGEOfVUzG36uOaY
4qH/CkDBzP7kzpC/KogAwt6RH1AoSXo1/WQ9uqPljtab/+wXlQFwnGEm9byRHZBG8/5VphnVascv
nUIyje0vyHu1Tll/H7I3U6K3iLOlZ72z3tlGFMdF4tiw2U5lRasJh+6c+nm5QISGOOhkC1KT7FMF
MXE9akBtH/Gaz3hC9VeARQfppKmLkz9a+87ojBsHtPUwKEf1nvSmaphKqCBTe6EREnxtScpYCcAE
K9ckM8YmNrQJ3jeuEt3Co698STSUpUi1lGKnl08IM5XHdAOkppUFvuw+++78mRHUsQ6eWUwVQxoJ
fIYGjA6v69lHb4V863RLtA+SzVQOWqL8GrNRm7cofUhyGrh3OvHxZ2L7ba6cgN5OElI3UEjsiGrF
yKue0DtcuAqLxAnQnBLpu76msOodTroB2MQf/KNA0od7lVJT7BnY0X75otFGM0nWoWrgKweWUdQA
9C4DesPhhp9z0nSPukFBy1a5HpSPhnn9tWFOK0b1Ol3Ry/zBVx52C2K1acT6w3VYRFyCZ4Uk6TCJ
ILdi0g1vx7vx950IpxwHxQOOD6sz2RZ3NWJFMyd2Uu/q44/KO5UfBhpV8N+AvHux+bUy4xkoMeBP
ca3lk+BvKj/l3i/e/9ZI5wznOVHRfRpdmNsIo5M1Oh+QTijgCqZRFVN+Mcv0c+he9jlb8kc1S1v+
5bB5jbbbRmu0YC57LON+xLKi5v9P6qdGY+ARD4dhQcuz899CdlrrJPtLLgK2uByucVQ6KBIsZrXK
tMnO+OEltpg7QUz3ENq9qtff7gqcMhISHcYLjpQvbPhULKRGHaQQ27vGiPdRd7hvNHi/c4dqjNgd
awZ7mbUtumMjCuVxmashwx8pO54W+qKBvyH99gI3rTv/D861fZpCpVBy+BFJMUeNbuGHF/FQRHo8
w6OjvAikUg3pEdINwEC6Lh2eMBR0b+cDN9eE8RB/jhnXiXE3U7JwK/Eqz8+CjTqAtLHdItA8ReR2
OIDMUvpGUW+hPl1ZcNfdWlvyQpchaEDosRt4HOr/QdTOYtjCMisao1W3UHzFPrCcYntAO8rLoIUr
q9PIOh9DP9DtSTiwHBFnNjlJJDCr3wOju8zTeLoI2Q9qvYa7ydNYo6M/CCsNLpZ511Cc8wJgRYAW
rfO3jP+9xON1DC9pbMUvUsE6CaBTFQHOpMJ1tnB1VrM5eHzC9XYKWq1yk+xtoO3+f9JBFrwl37CN
kg8lWo1ymlgbftQGk/tgZcZDheXMjvDykV8mpaq5i5s9d/HDS7xG8H/FNH+BzTLgQgT84hx8csK+
A4jw6zKs7tjuG7aEG25PKjyLJUDwcRLeU0UbLKxkzpydtKUJ3zfKuPXcEZp9Pj4dswmeGwyVGBpy
2em2khQ78Spsn3XRJeJyVNAcZaonEtyxX54drV7//YYgwCkZmEFMrmlE7eiJCqg6FQ5Wn1qSY8PD
2W1HvkMm30cMGyp/vj4ntuXVJv88FBVRmp2nhHgqyzqUWnAcKEkYM+DwPHnMy3bHLmCxIl6M5yJN
+lGDfd545+GahBZSobOq87wfboHXP/r7a4w1CKwMTZpGXspkK88rvHQbrPmr/As+50MOEtgfqC0C
5mWCWQpdEl40Sx16C6s3WqDPcR6XTJizJ8l/iY93F0Nu7bEeoALz6wIdHVhPl2ocdvdzyUTJA+ZD
dnskLMMgeSsMqXmxojQSwLW7HEdEkEexpo/DR2xDNUn+T6VsccmfKljCEicqPe1mbC7KVqgAjnus
lNnvkOT2wZUv5hx/KQtab8QPn7UN3kLUKwnQuhXV8DlMArMuVcqsfaKHvM9UaXzaTI1p6H997mmX
uXIDi4Em4htyD5TJ0IU8K/+JtHU8GqsOreQVKScZqq4zx529V2HQoMSYEXS8nc3QD1Rdyfg9R2et
X28fjcVoX4vCzhVNn1Z2Pw7YUgUm/D8n4zfb0k+SLlp6cTcG0uriZpJK/vdiP5Spjl16ZVlKTTIq
ZOGA+sTXZXrK3kC87OJOgYFbH/osce+lDWqcc99rO1LvHK3TVUGi145MPvnQrodqeVfomPSnu+1v
BF8caYxXn6hyahhEFasdGYut9+yKXOYI9RBC+Qc4qY5D+r1rffMDW71LP99TJQvhY94y79V5fZz8
68iqFOQuW2jNoo1hVH0nmCUa2gxy631+F466j8EW/4cG5qQ1TCYjZepQbgfhCzpFcfxVzs9Qg531
pfhQcTV7pYIisrYNynQEDCioIT4hIgDzmJFhhbMZHuxAJUYYVqBCFuvv+DcbJIhO2YueJ1z+Hxfx
vVie4Vi+Nx/Xopp1mFel4xEqMw2kltCbQ/rW9r+pvVz/vCHp8jCf9G3kx4CFyewJJWFLhGl9OTfS
JJrtnHf0uXIoRskek0SdJ+3z7YhpIPNsAPqsXISMwP4mZgnFgeCartxw7vyY5GMr2EMbc2JiscY9
lMWCjSzrIsSjGmlUyIj0Wnp/tKHt1IFnbADDmEBhUhwTxnmE7BGUyYmSU1eKLm7fSLH/AI2E+cOT
5tdiIt3BNOfRx5XJuJuQAngZ0C5nO0hb/1+irpDo2lGuNDfv6bHTIzXyKsbQRCNKeMyIAgDjKhW1
cTLKRH0WjBDcWiwn7AQ/B8EaGMa3s/9gXvQiOyOAKJ2vaYJtYr5M/vL/7V064ECjcCbYt4E+sI2a
CQN+vRZXxbbSBw0Y2Pr3hIa39VP/6LzUmxuU08aqAS0eMKEDKkOs6JRdbEMzLqrcDV38yjotAtfG
LtsrBqCEI+Tjb6HaYefvY9sZwQ8KH7CvhIm5xsgvwy6vzPyfugUzK10zKin/IDB74qdohVAmY7dP
3SWAtdoJ3yuTM4teyNaLEX7LuSWL8Ud4wMuQHBulvf+Lg1/tVyaI83kN1rvxb0qO16S3DpKORLsx
RoDI2jiUsnZDYSR9E66INpqZ1EO0i1zOhIdQn7bCHIJsAN2Tan2VwcO44FUmmmEyQ0QG6salCWP/
f+2R/pGyvR2cjFHXSQVMp3dQ/CBswrcexIAIy4idRqjP0r/4k/KkhmPQObFUlVe+gwV6Cbvogi+L
ojWyqwT5nBRXXBn9VqJ/my/jASDXtG6NqBQb0sDH3XReGI4l3Tow6C25DlvaC7vx4ugNUqy2IRk6
C9MRngi5AbG7v+aaNZDml4LwXB/cMzjZDF9ZpzG30oEoPPzala27fVP50R0KkTFbzENSw3FDFeNw
YhWLNKapK8c3IIHbk6HOLHarVyTmCrqhDHutyOhzF5Qw0tii4qdzGQcUTBYhpWD2g1xKVuCttJH8
2M7M6/1WsGIfHnQ9CYQTRLztfAVZowh0dZTr92RNb2MiWTrUeyywv5GHEoh6G3lTizSc6YLhlY+4
x1QjA9B6LUYFSGILzLmlQa1gO0sqEtcit2LbIm7xiU+5+F5/SR9e0IFnR2HdYjitXZ/IJmMeOgyC
HzMrtiPvZdC13P4si//oKHMiNLND4Un99H1WcPDQTddtzoGDLG7pgrRoKP+ZSCn7kH6XoKbgqCv0
/NWrM57r/LBi8z0vjGRIKsp4u2seePLy2A/WDx9+QFg30S5/CMfNhwBg7xxFQcCzYIvRKySvFsvp
n0R6S/rVG/MkOdPKPBnZQGwrOPZRi2+dSjD1tVhdUSlKAaEIesL+4/Pq6Trdal9zBfqGnkuknYwG
zH20GGbMthCieAJ1gO3VeKpra/Icl586mnZ+ZQrelwL9apnumUgUsOraQf5K/vgVZ+rUng2Vi9Wo
ByLbCfCAxh/K7A3N5dwutYU9Iv646JWxqWNXo6JIfqf5t381uNsaI6SkjrfHaYsOgof6AKLGFBty
DPqZd2zY88CQ2POyiW3SLtmMR3kt8P0czYmiTddnA19X3oWz7KPuJiL3SGZCVEqUFcZ8yJSMJMys
05yz96bS0syvPNCMnTlV4PbX0uYgg+kZ9i36w5amxlvdK/rE4nUiap9JqFe1in2XgtaLR1TQnDVs
y6VD5rWU09uWglCQh02le+HQM0YLNmyWWIP6q3r3nahvhJ/D4AigjcfbsrKnA3cxZ/FA5yOt4Hog
OXqLGPaRbabYYzR3mNiuui7DbxiUVgbJufvDoml0INjs357CDbA+a8UxHvqnI3Ec4Q4rEdS/8wFG
h6jT5pLY6igd2Tf38UzqbBYQnzOLxuCWLn9EHmdui0wA1exzdPUPLL8W43E4l1h3LzZ+n5zdwOPo
uboIe6xrWRqSNmTOvccEGAsW/+PKRIfUBSQSvXlTfe3D9Jby+dx5CD/ZMYWO9jYcKSIE2ox+U3ug
6wruyP4iUlyNhTlWTYwqzwYUQPmFzxsJsVmaiOONsvOFE5c0YISeUHpgwCLdcZOm5lpU1dCMAX/I
OTgN6QvkNcx9NLoMO0SKrvVUG6v/IWKXfOOiY8A2VO1NP5XUJ5aIvOO/xsyeeheew5nqDtftXsUB
HlLHV4kFYoBHlkKkgcbaFSiMFhNaIpuObfyXXPQtkcCVEMoHD00Vk+3DwZJrnhp/gWj1hKeR3y/t
+Z8juDX1GADg3u7O//TZMfnKmqijldFD0haJMwxoafw/8FUGbzOlpRmiU3itGqH3IBQFW10PFGHS
cwILqn5AWL5RyORXN54fSGytmo/Bgu3VzPjmps8CE25suJnk7GRQS15KB+M4E4dj4ixo+4H09WRZ
DaAa5Wy82IDEz7pyxUFz1LEPSGR+nPWbPZXmiUYBet23wKS+9qn5GjU1cTotuZqPWQwlFRAFaoXp
ZmvVtyaXC/7lhdI4/kaeJVg3uzs8TxNHVcayUvjWtRCpX8Dl6Xd3i0JNcVagJTyHcPz6vEadf00Q
2SbBBcjZt9gSbkEv8FAJk8BtAxlUOX9xiREEdWzljg7w/EVpURfek7EL8614NxRDPrpSbdeSjt9L
G4H98EGynbUDQMCrjJyxmZI5Z/iWc6hwagniAb6E2EcapVyfnOBJmenANSkNMaMSm+V8s3MM34Yt
xsRsmcIa+xRR8otWpV31OOo70g861kUeEvMwrQ6bOshRJbgDR54z5PUXqEb3H753kTg44DaZ90dC
7lEkMfvDY8Ba8hBKiFdL3+qO7aDBSSbpljNV6ObwnBHWH9wO92EpaBfzJrKb81lo5Vkw/sJMSOsh
90CSup+GxFZEH2pZfCEDT8YCYKLoUrtj+E8qVgMxgPfAgJD7UGVrA3GPDZ8zynaQfGBtbwg9ZkDD
rz4qt6CFhTh2/lJmKM4Q46rrWtrgAGhXudNxJd71nKbhTGqpE2swmyO8KggqhEl7XcMoId9HOnmd
cWjHDkIhylF+V4l7Zf6A87phT8U28gnhjQxqMz+t3YLQ/4CrzSqGoj0XwwDxqZL3V3+g15D04oVY
yxekELiaOvB99i/FqFGIsFxax8TiAd8k8ChE8bxiqzOnUyLkaKRbEIrCAaNzn1ZEt1xZVLBGwePK
ns5PPzkoi8g33TVhMRCkEAm27m7P8PQQpLNX8W8eXgPbBbPRaneWKRtfz938L6eRq1E9ZEmCAys2
iuwIY0QmqhHITx67Lo6uUOWiMDBvQbPtEz+Xg+xc4C5KMkncWZQbD484PJSHH+ytFfrw21C1zle1
t3gYU8Wc0AdkT4iAzDDqPzWgPjNuxKWxxKoWvF8Y7Jxqr/PY3cKqZmpIJoDTNl7C25YEVWo8YkIT
vcvDTMPDkSMl8WUvrn1vnGZm5cDCM1OiHLdpHwsvtOl4wzv0LKjQxODmoI1JaWyQjZD7Z4WL5B2e
8gfv75bR7VPkZa+jfEZhHi+Pcly6ooBgxcSeMHMb/XssaNHFUvqEh6c8x26kDP4SQo4GqFVtGEbX
YSUwR1OByN+whj0IpXoHM5Se9sUmRzAxs9kGRTK9JgI9lGYZ0mSH34D+p8rVlf4vgOdfIUIS2b0S
+mIudjqd+1NHvgyybt1K/O5pZ4GCChvJIYA1nahWY2BfcxY0mq7HFMKbAiAqpCVcL91z/odXR+FV
41sDNI0DlH14B2HmQaYAuiFXnYvytgkZ29GFPuWVExzZUxYEuM0Cnuiq5kw0+jXKiiK8oIdgNyoF
0or1bcfhn9/+of9r78xh6bcdhaxO2rBlMgsccLX8D1OvoG++Dt3LYmQ1++IoprC6j33JIa+fhIpQ
bQCtAh5JnLzorb+EG0fRweZtmuiafK10nSEgfaH3hsP47SgNTaNpbxw0KmkVlYtOY4XPLXn8k84l
VGMWxH3W8F5DZ7ImoB/IXmFwrSQabI9XdomjzwknVXCU0TjiUXvgnInV+aFhAAfMFki00CcjvW9r
gnEj4r4dXapC5S+eQHilbWcnH2FpLeKx+zd7mD+dtmP3uxMY/14HrwoEoh8SYvpXxF0xKpshA5OX
pNP4psXRps+mbqqGlAoufvhN6gJyi4o4C3PyhNGpJIXF25R2LZh1+O/auLPiYu4JoQ0w2Zqs/37Q
kHFUdWGHxnElG28ufGGJ8O1ZxSb2kkey2hieiyYH3lfpDqDul5FXx1n0JB0GwctIDNzy90wrplTJ
LlIasMsqty+PGGTNQ65v0eVtV6PEIze4T6MYnkGsjYMI+CCj9JbzSkIuq1ODGuLanJgwT2SG7/Tf
pPzEfb1EauslHCjgUlC32Pm9lf3HBmObHK0aPRiTCdISw59acLeadXMBPPiOya8EvyK1ekDPwRRn
Jf6wIskBDcGT7Rvp3cblFp+eLEjjWvH9VKVbWj6S+NXm9PlGJxsFLRzPenkLqygocIsAbA6zUhnQ
Jsy0edTONiytsIMAvNfwKPpb07DJLIthsAl5zINUhPGWB8H+9Iia3WN7o510PDpWoQEuFEN6XMIE
k29skY0vlDSNm8U4jE5JTiklwL+gYsxmMP7iL930ywuTMHHRdp/7X1lf9wHUm/rInbF82TqXADfe
xenqBTT2z+aOkmZOSMweSgRWYlLLn2aZ6UykajI5FOM+eMMy8925XwmVAzks6LGiaQ81zFUYWZxF
M/s/U1xpIOjkxsmKDaW0wFN6pRibekxQaXxyOD0Aqbw0EmybVdxUpPjNxE82saC9Wi0lecIHcHhE
uYWprfB9LvnCvh6Sg3Nfh4SpoZClESfrTO/5X0Qq7niupPO204hLxEeFXahdpllNtxos9F6TSyO5
UbHaAYwOk1vyaoUsHQ7bsei0IvJBxAD0H9RP+012Pglz67HApiq26zjwlv0tMfHLCHrDZv6tGlEm
d9fgSYh4FVPC7wJV48/fq27B4z9YRIeog6MgnHc8Vnhha5St6WV7QzJyh+WZWjD55AwOlXd4/GLo
76CsAmRnurQFQwd5rKETFIPuyXTkR7bzl7hKq/eYIRveU5xVLEsdoI+jntMzoCBm8khWFTE3ZMml
KwMr788bvMEqxhMkoPfuohb+HfYj7TFQ8Yg15zElejFgz0CMGyG5T2kr+LdnquQ8nzbw8Hi8qlFX
bIZX0uC+RhqZuX7019oyUI1q4xRUwSwwZikkDhsYpDTD4kh7gxNfLXKQYwKOj1GoWSUklIYgJ5hU
iTOI8y8QjBL4TDY5yERJjNoBSS+Ho2T6DHgF/XD05SwNQ0RQeZEWmBoPTHLpbSZbSpKd3bYg47GR
DhSHRiOmgTPVvbIJB/ni+eB98eggOddFFP5mANKzIkRUtBws6TyW04bcukHSI7n1gLZqc+neoWzQ
n0tzECy88xRBBrCF8vbm+I85CEeGMXKVBvgLHptj6JSOcNpKCAT8Mt9KeNfjMjV6guq4HR/fJPFM
LxhssfJvz1CyXsSGCH5VbSpYXWgVc7xYVTuOTNxQcGVpHcjMZkZfKGJnyFBeoYrwpPdEFZlETUUf
mscE+tXx23EnWKHqpmq00MnQKeH0zhuzMEwf3eRdb25ksDwaZQqt/JwAhvtgyw55o2A1O/xTjB8P
kwJAOQkp3bKozCNTbGM2JVY81sVsd2AOXSwdKEYuy+Ebg4fMv9hINtjxv9gSfN5BUJlW5uIXBR1p
EXbjOvaJksW81p1Dg9B//qtF2W5C6kfAgVIxqhpq9NsLZoL5wP40PM3tPDwcjunakITWBS5k+wpV
jgp79z6+TFOFSc4LNI4u3d+AlhUpQyKQfyeCIWL9lzcQ4PeGlSFSIwHtvLQQtW1+7ZpgnrEg/sOS
KSDFXhKHsvsX9HTPscwsAcLeqVvYnRfYeANC9tHgvTudWfaetCAVgXNKZa8ZOBBJpEGVCXRpyQyK
6u6x3L2LE1R30ko0sD8QAlAu5WcNxd7ZwrPsFut/XsAzf+xE3UTqSJ442tXq9yuFE9apq/Owu/l+
/m0KvhgQaoqFKdKHhQK403WxJk5kX/6r4+KegMiIXBxbp2AcQg4g1GWunFy4x0+QDDUEjR9jyhbB
39pdrkufxYdjhUYfzDpngk2yvutDzsk4kETWmHfQQIwaVsAgFUIwcNi6rMl7avAUd+94pumNAyD2
T9+FS5jv5yhGl7LzZOQzX0znqW0sYr/aQcjm+F3IwkcxpF8Etg72bgf1sSEBn+2G6vv32EDiGzXa
bPraHjjSPu49ri1x3vMLgTgsWx/CNw8yHrS1gwQFKGMm6wbDPVbwcuCC5lBvPkiRu6fohkyK52VT
RIA4tfRZ+SWI4K26tGzJcRZI3GQ8Nsj1UFZ5QRX2Z9ZrGdbL7CPzMuuwiVg98ttfqgNRY3sz3Cdr
/oufWa5/tPphdilTD2IvpkqPprYPuxAggI0s7SduZCjAOvFznYrfaGdc+oMNZt+nkZZS2KfvzGc9
rB8AeBcnZXi4D2+jMdcfjT9G5/M8WuUTlQ4f+btlasEB0gDDLwzF5zcfyBn8e5m3pcv0dTXkKX9S
zqg41rBcF77SELx7dt43x9OCvd/oMmjqXJyv//h5GGHO6WXU3PjKYR8jiyFDaSAWY01R4pat6xf2
GDOlRTOjOpWY/QBY2oCC4y+e1kCloum66dSk9g01XYZ7XQLlPHVBSVFywMBNO7+Yp/rsu6+b6JyE
Ozxl7eHa9zGHErELH32UAfk05sgNlmd5kWHBdCKzdCC6bgoVZvR37bEf4ZiQr6GrKG880XxrNWhs
YphvamoBg/JbYMeDoAKzu6GgqE/4abE+7go6WoJv/DYSiXOXiAfx2U57hbDLYywHEMBxffQBg4uI
lYLVQpYU4FBYQScTFfRIz/T47rusOpHHboAq6pBftKjLyDzE1BJuGg5XR+ndxxuYY6Ia+u3i2YlQ
g50pG0xiqLW3qVuprbuPYpInTtL22qSRTArO9KwAkFPx9rpS8I3NS1nboo/GeCCXoboiJbcDsOBM
cyor09xTQfkl8INjZLyaj5aiGFvCAEaYhxyuMt3b+JPRB+MPldtwq1Uvw8/YDtUH7ge8Pf652UUS
E4zEY5D2ci5H57fbBvGm3HPyKfP/K0utR/20ysu2+WYXPbeHMzNFmfvZj0fJElW/SSp8QrmgCdDL
FbI/qTtMekGq1OXwlK4o6UysNuRB83qj4aAsuApR2YObNUDlw5Bz2FUn3V5D2tx51Ke8Y8pYVlPk
9YIaE4fE0q5UTOzHUpjLKjn6okp7YcBlHQicoVJ2rI2QCZSTJkHJUtm3IqyLQYSqkjaKRfPpp/tt
MmP7DzlhKBTuHoMd2T5yvkq76ceTM7bK3KSnEM/KQMGfUZ+C3QDsKydra32/TUrocyf+eKnvFps4
H7DF7ZB4rNq4jLcHmVomrkNOtsFnIYbf2+PNETRYjWjNMpn0eDhCSHTLjn+XfAz9jMaqwhplG3Ca
Zl3dJkvoZ+7UX+4xvb69oKPkFGzwWRF5fsJP8r/KfOagosMAYlS0wgSmLiArEZDTomBl6d0I4da/
JtogAKjNVn5q7Su76Zhf4NnfDivPQlX71x+vEqYNcK5MVvlp1ej29TZ1itQ52TOfvprQGYekf1mQ
KsZPpY501G2am92HJPH6WoPi3Vs3Dec0/d3lzPfI1szGfjgyYk37bfQdX8oPZKjlwxRtdDTyQhfj
GACgD7+J/qHt800zJztJ+BEai9mU4o9fuyEBzw+F7vXm8zEwhgiVZzZQhGgaiKvYvEvJKsBmmS++
ayuZ8mYbbJ+Kqhm66y4aLjDHGPNxFPn71QJlhTQ8LapzRuiCEZa4A9N8Lw2yyCLpbWpHOBSDYnfO
2WWKBdptL5nuKoXwXB4aeb3M3uH+WRZxb/CS6xKMpIHuiJ+pHKSx8JvrGbn/r14yDwYxjhbPe30O
9kSHyh8z4KgLaq0pp+qOol4TRXM5zv5GE87CgjzigG9uVTnezFRY7P5moHwof9eJqro/h1Z6Hr7a
W9QLwj5dMp1VpF7bL0JXN2doa/nxUOhvvUfBwsGKR6RmLciD3O5f538efEnNMLRCD0cWgZgidl1c
eXLAgGiQSYY5OhzFsO+Sea+ee5P+n7MVSY5dNwdLgCVNu6I0iTDeSaaSPfpmMet31w+5guvj4m80
K+NKF0SBCGsEgGGWtUOjnuZ3G+4MRMod6SypR2kgRIeAZepMjl3GtOtVThgnQjmUMfPwmgP2Qkee
ZcZRBNjqurv6rQfQKLIZNaJLRNRaEG+ut/ZZ4IjDotvtfJagagB1nEBxgX3jPq7/ViLxKLaCAdX7
MR7emlqlWl0VSGDy3WYWnzeqzZNC5dcQaFtAj7Frj2XYEBupqg2uVkIfTBOM+P1y4PkdA9Bt4l6H
x3AnfsM7LRo+8XQaBxFvEdbPOe31ohFJZLzr+ewv5yRI479ahUmI/EWEDiKEKw47d8YhgpqMFrqF
x/9fdIjPO7Ei/2WfpA104XUxRN5GXJkX8bBt6u783EMCXGOSmEV0imeVkn0OxozJ+uhNy+gt9UWi
gkSwKflORk1PPpSYH5ZpdVai7ESQixHguAXRkztFaI8Evxo6qCieKBgSWf5VfHN2YSmhuxMqNF7g
eWYCuY7z6Smq9qYJ0Irkhdk9P1z0RR07QLkt0jIx9CCfMYMRGl5zToLPsn3s3PTtWQDfBoc7Y1O8
HssTB2nzAEipM4iKYNKebDIAsaS6AFf0kvxzzYMCTaxwU/FY4ISjZuzVVTzMNp18nzH7Ti3P9hXL
7GhYsavoiuMZbNFM5f3UuwZbgKx/XXcV+19ysdZTI673xKCb2R5ArbXBMETAfIaVbax7i1uc+Nri
TrH3jvyXMax4E4zzHK+ttktJ9J9H9ofgoh6OHp2zdL2zOQ7yh/c2QmLxGlL+q850Y0K4qVUVA9sY
9H2P1KT1vkxTZfozH5n45MLFyPXTRgj/+sy2yxUM02gPePOcrJhkWelR45x1nsPp2Vb6u+ChS8uZ
/789hrzcBaPcpUy+4AyCRqLHqVVvyp4P8vu9QwVHDPlOrrdl5RItroC7l2Tvmp8QPRUMc/z2fyXa
ZyqT51XQcsKVDreagCxnh9FTP1oneUPDR/Xq8+7aKTlY0jtKWZKrh9yVAr11M8TxFBeZljDUg+I0
LJbbTdq9CSg9uznCOlJuIk58RJLMGLltkV9kn3pmIoSj97K6/1xBPUIYWCegctedToEIzM8HEmNQ
F0FeTRh1emMXyQ98QOr+STH9YpVUyaLOsXhg+9+wsOH7Uht8tvz63tlhJm4hVwvZ1UyRrnXy7+el
sd1VawVWlRZ+BFPSn+smPERPJwmNtBekHGwkM1bTWQHTEzYjN5DsojC70eYEzBEgU0RGjk1l6Z8i
ozewUBjyjoi0Y0zywhyCnPxSNqtK4wBuNUjr8moJVuo0DCp9pTgQqB6UEpcl7nzKRcPSrSJjczBl
9Z7wVm8d/NQe2YTELrPT+obrX53gLy1JU4FuXTI3iDDixacMWRVzwIdwSPgWXhGlCqmH16Hvse40
sFzSMUolV9J6+w9WIIgzgXcyHlSZu1T7OSeEw+IQH7EwyPSC1yqWi3xKfX05ZqtkCmHDqVsw0Hpd
TMw3JDqNqkjsDF0luA3CJlZR10V06Rsb+tQKd1Oo2pl50KYw8NTd9LP4xZglLNGroz8tqXSrgxs8
fbjfH/zGKPFK1yhK+4wGyTmbR9yCPO2UIrhWykkSGCWpKFViGbnfC5wXtu/2jsBtBcKTsgKLFrKK
cEpmeF3FXUCWqcTzhXn024Bqj5wCeVwIu8UVXucvCtNaJpYNezgFgFXxGkZtDFp2NEo1QtmSwj3m
dnH4RuDIkkOfIBDg+yFYxUc6VAlONPYJdS2Sbut6/eLc3cdS56USnTTkZk65pY/bykE5atkHta19
I002YprpwWi484J7ctkbg50r00UxyY4F1KoLDDgtLbmX1TMT6i5XpkkZrj4iwWGA3ZD83xP1osBd
RKvnZ/SQQzQGra+fUrTc8pOUCZyYbiSExXfPAs8CHFRx98b3EQiMi0AnJkOFGT5XYgkAeSyMpbwR
UEDzmOCaDXFg9jooDdZcz1YUZ2yUn9mQdyjUfRTglxc+HBqP/H0gStwH4mw8o0P1pf9KJYmaGC3p
AqVmBLNARO57x9JkRESEbiozmoNVra5GURI9da3MgZXbyUrnpbDCE7DmGduWbSi1iDMb+IiSKNpd
lOMNEHdyBLdCMJNfI+WE+SvWU1zTafM7Fdig7m5PKrdbodZMAWlNUeujG/HcqmX5M1uqYzDNLKKM
l0+nwrqS52w83Uf/orVm5KM+ECyLbtqk7z4Rkbz4eamJjPfFOejvVszpEB02+5VBao9P3w1wuVAV
JsTDeMEU55V7NrJkAcEHy5Ycy+B2VVHKLIVAyWameQ17aVtqyCBAxT2d6uhl5gObZKicYHGt7SWw
5S9YC/oAGu6ihIl5slasfu/XkS9OM4I3iPsOQNcv3IiagP7BugvgSnYTV915qw6zIT9pJ0mvizuK
tE9eWj0GAHwLC0GmjJSor7az8eE12+iD1IiT1/axmGV5G70OgMWBlOtvCd1Ln023zU/X6LHGWs7J
KZqebo20HXUHvEWEsCh9asWCvV5pLUyC4tSK2rd6QuyhE082/s4z2iFBI4Q6dVdEJc8zHrCDzmoN
9RLUtEX7h4X8rUo02/CVMBECYI/dFCSFNbNuBU6NXaJxzR1geA5GmjAmlDstgsa47cUKHDcLU1Gh
Q9ZYDH4/rhYJ/ljRMdEOBRwFTAZhDVDf7ISjbImFZFAUupPXYPUnEXA8zHme2t8d4rjEzipDHQYg
5F97hXvpKTFDsskRmeXKoni0vZBPGJofuiLp9siAbwKa4MR4CY8o/Imy0KcFeUC8oHHEswLfxch7
MmsjxbrgraRepU4vOX9Yx6MuWG8VN2sxaZtfpdCZSQ60B4OwGlrovXKKS9X9ySZfv/Ggxyer9c4g
v2NczhAeAz8KQ6OJ7z++dTVbzJ90bdwtWih5HcBsui6ysiStqauMgrUHapdooseDTRvBcT/rcIZ3
ye4IclEvUUwNx94GrlnIGaW9104YL7JxX0oAIQY4SHigQc5FFrqoz17y5S34JR4DgMUabV1yLa2t
F6SRI6a5a/V7hBqXZwUrj9xR1mcbcRTNIwVmg5WZqNKSyINaSrg/yr+mYKw7rNkuQYgt+ECvKnmv
DFVpB9otK1xq/qQWADrcX98BIcxj7s4cAizJIMQW9y7FCXH4aNCcZ2qNbO3rhq6GDVycgGqZAYSO
VOqXTcpAdb/gSnTGKfBl2XQPIRtAOKMFKwkmyygyZvHMMGAeZXtMey26nd+3wBT7URfPfgUd2IaH
8S5Flmr7XArKkI23+c/msHd4pdOe91ESvr9CA1pfU7AHQWW1vPt80S5ajsbQFACO0oWS79NZNtV9
dF9gQKjZlX/UixuL4xjMB3B1m1S4/DZZsEpGXAy0+8FYy/G6zvmD5nBn1d7IsaTxQ1sneDqXGaKs
aGuUE3c8BXUXSz2G3IoD+nMjD7Wr7wfBzt3Ze7LceXu5b3Z41Dw4bXAnlau9xKHnFep83Yt8afkU
EoAU/reCtJa6d8S/PjTCwKSPpWyXIV9lRntcIFAOa2j0zagbZbA95DGlmPQuCJyOjbqMOb7+DjLn
KphK5Sh45f+uAbsyF0tDfZI7ytFlI1h+NFtx/WV3n8bY6a5Zb/agoSyz6DSEwexLfWzeZVizfTei
Varl6MxW5HRHJG2/KHBvHAMGB/OUbfu4fsriwoMgbmO+EvzC8eaT6CVzMPFXMdFGpc9BA339rIxs
COTPZheDtoBBDmDiUXpENeSF5fnUvGDPAvKrNHXBZOlMgIye5GCYlMb4ksd7rLyFElNZJ9pJ4pxc
QUeY5O8SRzA+bAFztP6IH6lCYBQ1ey1zqaa3GfCTI2heVyeg6t/6lAO1mle3UAKXrCsbh/qlvLwO
nOg5OTSz2CsaV8S113+pumKI+BFJcd8g7yXWCRhSVdMPb3S1RosIkjda5VeEA48u13l9ISAEYqll
asNgUwTn8tShfFcC7IpiDsaytLroTqf7uxzal5Q7myC8x4AiQf03gcvtWzImO/re+P5Uw/FK9Wq9
Bsowmun9lou+J/7u65L4QPmMc/Fey4M6Ipou+c5WSrYMNSsb4/NR4sE8hzpKUc8s6kTxPqg07xpO
3AW1xsGbU2/KK+dEjQLg9r68Sts9gKIxZSWt912gIFzgWOJjZwbHvwn376xJ7Ngjp7Nue3PVJRna
3Slgtpvs8WI6tvqQGqIFZSiZIJnb8ZrK8qTqflrx1a20dkPkLfUWath+9b9eQbvDkFubBbJxpdqW
zQ8xg2lARMjXCymJstcyYGUAL5s3HfZT6NlWWkO9vGhnph4zilO0jA/NCjWlaYDLYyrkdNPK3Ofp
jpI3U2VeRbwjRUR4lRIne0OyohphgQJnh422cLoWxY6nysb6rwMXBAMCAJLOXMiGNtZIctYZUkzy
Obj8na/z31dY/IWvAaDFkRiu3KpMKbNhRndRHHf9T/A+95Ri3KY8aeP9LOfOKQkuXGPtwQlBkeIJ
+BlkEHsuSy3m+xR1OPEyKB5Bx4un4SCoyXFpxG3Yy9/9eP2RCpfL+PT4O84A6+MfK5XYr2o5nzqG
5bkI8lI+T9Q8G+f/u/X2PyxugtnfBLlDTPq9zHHS64tEq4YO8O76Xl5F2K/yW4q0dTZ72qhGAlIT
E4hJnTrySA3YVr07gRNXc6DGjm2R8rqu/Smv9etrs5+P7bUnviDi+OoAMqaoN3KA15S0vUJUZe6m
CUsC27TY1mNHVp5pZqK8rAF5IEoyjDy1DAb7T/Te6DmLEPSRRP+1sqh5KinGd3PzdSf81WAZAILn
smzLcAk3JMJ25I2J2CQdCEkuTSw7O82mWxVVVnKmmpLHoAM11ABRe6Kt38v59vbEWAM7ZLV3Grky
6axudvWziiSnZbse+UX2Vf798oANgQFRe/5ba2D4Tg3x1pq9CXy8s1sxINgky/eq1RYCAZEs2sAH
Va6A6+4PWS8+1PImktKC0yq6rO6o7idEksURAj1AU79IiwSnP5F0nCBtQfFfMROfvJnQ21nTRzcx
I5cf9Vz0pV6NG/YJrMipgT3IB/vTDadywugM3QqjaiiBprgku/7u1azFlom7myNkeHJI1L5y3i6f
iUEisNAu7DEDdGdDjRxqdtH/J7Pp7VD3B0KENspTEG860DjSvq607XCHYIHR5tvpaE5IiRwRhhZO
MEoYsGxQSGrTUxurSFdkO2+5a6h1nCGeUHITH90a7rvlqhg4a4IOJkzIUadBNoDTHpAda22jp6Pl
Z9Lxi4fwY9BNrLItJd+wFFLOBinl4K6RucS51IMghg66UK8ZHkwWn0qh0FiOO0VvZV7wE5Uhq4mW
X6CTJ66nYNb2yyEKBX5Az54VkRTRoNy9FCmAYsJjkC4tpz7TQdQJudHX28PBxQnMAUsN1lnYsEtl
n0Lrcj/twMnVoEzdAymZ3WJHtvFyhnZ2wP0nDhA7zk9KbtY2VwIdaJT+HaDtoT5Gb9tTFcVULIOw
ZmpxEJGpd0GIg9GPEJ4kc0b/0v91/JD5+JjzYctfQWRptA68S58XePuhnlgzaUsl2NvlVqgYY09j
vNPSE5qxF2nSlxMmutRsRVah+MhIAT0ybXJQOx2RuOIJ2SbFZpIOA8LHxSMbTf3yZddNcwXicGSS
9wnihtUS+sy+9kJ6cvfzK9pE0Lhb0Txw9X7KQKGqKDH9fBgmPbCHkJH1qBhmbnGjJCveBvv9BQZn
VfEoMSPPikHL7KoayzSm/Pm/LcPflLtQsyeiymFoQ9aH5W1hfFLRBj7d6gMermJD4lMnRTnXBMDK
OdHh+pFDkynbHeoMsZeQsMNrZL9H8gOI0bttoTRUv51dywpo84EVLfLF3+0e6k2SIOosHiZnkHgt
Vnd+7FoHK5K+egWEEwyXUbdApVSg55EIFQjls4edXSjLgliwLvswoIajiCbh0VWyFiImjJ0/3BlF
W1u3XcrXx6m3wsHpmT6tpdGBsrftOG3tlPlk71q6MPafN/bWIjG1waYJC+5Tfgp3cnlua3DLqyDQ
xYusd5ViOcslMBdwD3XOWotxgK8ZM5HMrilWXDFln9hieKnmvK0zs8usQOe0jY8UdDlDgQvdcQZA
z38FwX6e2i2+SJt7xw8Zl62hTql2Qv/1nAGopsMuUT4Ry5kwb1+Ar4o73sbF8+CrcZvkOhfENZ2m
8OqjDelylX+ogfN3aLL7lyQAvR/Xg81xEDKFMlzliRxnuJWZBmDo7Yh5apMAt1S6grUccjrL/Jmc
1ytUqK8AV2a9peb0PpO3kxy2OAwpqDLIqLoMy72jIvMp8vIUh6Te+7QMi5WNdkWhi6JBxPnjjfC/
32XeRGjiqP9+awqmHQdIjz0invbwEyQmwOkM3sm/R3oTjwYwPs4iPM8qZfpsJzUrgw13nTq9oq6j
xE2+Ynt8GnRfN1ALVVwIryePF4evqham7f+mj5Q+Buhz0eFwsG8Mkw6WlXP48uFmZjbzYHGW+FjR
95XubLmcmpGnJz6FKEUbNZV0qZ6yva2JGEpFZmU7jFVwqbq1wLScWvuzYjL62XYqDaGq9pDn8H+d
i2oVgHao2TxCpeGaLfbZhX6L0lHQ9pLdbmo5cy/i3kinA44rshuyJzRvgUgoQ1m3QYa56bNWphBj
vGrq7woj2382PqD4IwyPYRENYsa1LRKBeiY42B6FgKzuj1qQTyphxz0OjZUc4Rk1ghBFefmkre0P
TnJ9RLHIgOEKbOw1Zm6C6iI3CEEHUcvE7xVvLvV7gd9xYyaMMeikM7rlRUuOgmbm7yWRf2Z67qLv
jzcz1Hp1xs24KncOkdnp73FSkIFBR833bh8C216m8F6TeTs9+/FQM3/fuKSYIOiUDqj9VVH162if
fDwaV7/tJD5MEkYkO/gCyXxHmkaMVthox+m9+FfnR4XkQeq8in9+9KYQE6aq/Y8R6QRaW35bEwiC
IyyufDfa1Q2dT+J4raADBziyyXHuqbyjelY3EuzQ1I0GbVrtITSaiJlDiDD7TftfgPLduCRu/93j
e5FKZdNcxBD5yTC5vmiXdmOYMsBHIh9l6GBTRG9zb6+39prNF4oG2X8mluZ9qutFILmifXzCgoA/
Ipkq09M83dkxHP9iuUhPqCn2Q+IbJvHRp8PaP+yU5xUJ6Xo2mucAV1kt1zw/s+15fLaEZmEeYy/C
PgtHBIKPce1AL2SwNO5/HcdgsKCcwhoc66VPatEi4efHrGlYMF6I29aSeJ/aVB5wPuo8e/Ufzk5W
eQQmwwFtBaxy3eXCzRNzzj6c5XhaT67MCPRbcRVWnkq2sjjj8XMsH7T4TcActlbIKVkvI2qZqGAN
MUGcUIR5qRRn6stPga8rNe7DSBx4LxNWD1YQU4hIP/PRLH7PEOXkaQdQ/o2vD8xss4Ab2KRajVZy
3PAbrboXQ7CgixqVfI5nkzlc6e+nXEaSPseFcgORXVn/I3cxw0OSt8Tyrqs8unF5ri4ixs8rBHtD
HyDA/y3y9GEgZSIRFZ+5UOsJjXs6uBXz4wzsPsWXNoVWfrwaCwOiWZJVhIDTyyyFbIptoXEEAIcn
nWU5710YKXpJtLwk9f+9XNNgrPyOZRV8kClitJN+0vC4tPmR1Gok4kPDngGSK5smaJSob2F5ZNyc
+4xrrmfc1WKiQa9lU6zsgwgM+uyKDHqf8DviZ+FE39lzPZkMUC+3Y3BmGlEAkRYEhv2IgoLgp+YY
BqerKHzgysGm+e/v9Hj9Vm0pHzmQvo04bhFE5ApyJZoFxm6Ok/nwOUzesIkqzkH452FxSCjvO6KV
5c6vtQSJkQwzySsCqXRxGa5bYSU301TVlw1nRa15ALt1Xfc152rd9mL2bAsWdpow2WrivUtrlKCM
qa4eF66PWO5lFKyUkRbmV5yrOS7Tgv9aX+icO08jTTEcSSruQEzDhF52XaFuIADQ5PaTDMgta+Y/
P3A3XiLazSD7HR1Tmxv3rwiNFBgXQDE4GMoGpCmjyabmgA5pR5ymnfkejbt5u0soBZgcOagO4tAf
o4AsHrFkvEuUTR0y7BQb6UOPSPtbJGuwQMQuxpx1GuM50kJ+mXN6oY0QemiF5nA95xrzOiITFGmD
9U0VSg69VDR5oLs/PUAByj+PKtJ1FcRoasQIx6lOKX0sHhJKi/h0B0LbeBG5cMcQMtbNnnWi5LuB
/cNf4s972lQya48jTubQ+u4Fs/Mvk8cx+39890KF4RPV4gXC2Qfeto1uCFxXhxY/2CmAhzu0xm/H
jSl0j0jVieRAIEyqZ0WyUaBrGb6TfQhlXyY9l9GlzhjAaEmZZyEbhp04BIiQP21KWjuu3UXkhsFg
KTOR1eVkX08qCr1FpnLYAVEm3SZsKFGMrfNw+/NRXi5E21tefV7RWaL50Sf9XVEiBzpa4yqilts8
YAMo/8qBLYSFEMuBqOSDQZfUL4mn70n4NSJdpPyMlsQ3M3HRutvuvcVWdSqWVzX2RFK7xl+NWhYT
bkKV7F3VyV0VlMbeQXF6vSbSbESKvGdQtdDak0L4H/s2Zm5z5K9a/GsTmMvakLaiGdh4ERayxRY1
xo34so0BzkLmB7mej0+BDuCKq72RCKGtRpetflKOiF7txB5wEyrT87POwdw1iVa3Qw1/XLB7TWhy
joAGxqX5v5/0rx5YxKdDsXil3TzXyo//6T91+Wusv8cHZYKklSporEMl9LWEEiXpELiY/hgGOyg1
1Q5VwOq8Aqfa597yS/JOkG2XdZIdGFdFksilzv2UWjgnqLQ4ZtRVs2/+TNm06tbpl/0Fhww/4ppf
NvxBJPSXm65OOodeUmJDnzRP08nJEjSKTyBxt6WvLdFGVS2HrMuR2qvMwWlxta8XJ/av4+lc2GTy
umb9FXwJpJRKObzfpyN4dWpLAPBsEIpMKl2aOJrjomNsxd1Txhu8EPh4wltnj7tELNUXTqoLP1Rg
erKcXaqYllSMH0o3rZ/ae2NtrzKXaqdyv5vQSJfsL+/voUpJWruDLPBuSVGM11fO4Z8j5aqEqFif
ob4hUkvCw9U5Ga5VSPEJHPbeQOXgbtsGNoqvoJaD9XVHMK7MzNJrCsnSrwfxXbC2Ul036WjpXJp6
IE0HE9xx8N8UC/elXaiaKzITxOwt6WflBB5gmBz224/COKuM2L63z+HhO2dijfRCbTe0H1fj2OEk
JkSGN5+onmo8G6LG4HLE0z9ZPeV8t7m/zKqMPPfNVNYS0zDNGHG56j5HLRHuMI/cEqhpYIU8dT1Y
gwvicmANr3rf5R4JksbNUhbT1oGMQhLjnqRE81iwESqhjvjWB3rQu3Xf4imGCJWKwFINmenbmwVi
sEeASHD+g+mpKpVC+lV+B7cNK1c+Gd+u4qqeam4wpPN4JcMrb41G0AYHvIpBABxxVPsr4NXz+Ts4
wkcXE/5zEVCQJheT2kuyC4WHUXbcPjiO27hegQnZzP1RsTbkBQl0NFQupfz2ji8HNFQMcwBn1z6K
tLl0E//sowao9r7wVWe2SvWACrbCpcO9nGSzG62zZfQf1PgSSYMF7caaGu8ECLxQFqjz5OmmqGtp
cSU/GGu2Xu9+F8/meO1lFCklEQmeb4Ti2higkuJvUKie7AQS7HLjG4NDUH2JG0Rmq9Xeqazt4/LM
4W1iviwF+75g5qJ/K1EAkM5l5ihrUlKLy4se9VW56QP/FgbeeBT0iqXexz12kznUziYSRaBgnrEg
5e48nMQY3dpVl1EpKLLemFNi3i5BgpE0KUmoQics7xAiSzLvlpCQeryWuPNASM+UYL94hbM8ivqW
97shHzrTDbMYb5dW6taJn3u/f2uAN5alUKFrVFDqBq9XXSXS6LUSKJ5lAbn6qfiEJJ+2kQfrxacx
Wk8yb4xirl66DWB+Iu5x2WCigul84Yr1QkU9V5s3ljRXSU0tni8RPOwRel40tn6yjrN7MLxMFcl9
CMWdSCGheiQ7rxljsFvTQ0jofH6VoER/2NvPVMF4sU6n6B536OCEGJcygoEqSDr4H0YEwt4eO3vY
u2/op6I3HoYVRaN1eHjRMpdN5yS6WJx8nfNxVBx7c+obiALuWQW6akLn33BI6/eKvFGopUFp0cnb
4U6zmOW+i6XkzdFYVQrfJtxZuCQILP3cpcBe5qIoIrURKbNtHQO8scUaDzIs25RFPRybO4WQxkv3
+RNzW3obenDgh6qVF9BFsQWdcDcJKo52S9uvjwoqOFQMd1rM8nDESCwzsctAMIQZDQbKnuL1riMr
Op3sBWb1RSG2eMRatrlZ0U0nrAqNsOZF2B1xGlfJ3io4FySlXiyz1ii3DhEMCmqDjeQ2ryTlXvyI
dOut3lEo5pQFYziSw+zkmB1eCVqm1+oi+cgYvSRKnoTVvR0QJbkLy9yELZkr+xAoX1Bn5zEaSZ7E
jvnuGsJCpfYmXqVWgzSC62mijIyEjRs9y9HkALK0APZ/b7rLFY+eOWYqUOgVT/rnUZz3YSPJsHZY
kwGhBx73ISZ262q0629wJLzfFC2krFRfLizvp0dGkMp0LD2KuknjRY4vA002uF1pJ0I258L2O+XA
GUKNq0yrSF0inWjOfubEuZOZnn6hJ7Q6gFSMgk4yicTMbIlD8PhR56U5EMbkU8Gfb+gWWAfEMcF4
3jVeykmP72S+lR35g9gjjITlcrgw5IxgAKeQUEf3E1xe18LQ8ruOXb2PnwMZmdW25A0+YgH0AsD/
xwVTvk1adVjRv/DRbiYpqg6LNmYJ9L80ZvtCuWKHkzNWEY+UU7XkxZIsiuZ+7VWgNkubWw/0Atns
CYZhbWv6atUZoi3nQFVMK58kQ3ZTfIOJ4D94p0ng620jjcRIDsyredfOeL0c7/fYpUyqhlrcByx2
aaC/RFtBYXcvztBtp272rIp1PNbwIdZ1ngKqiDjobFLbTu2y8if8G52dCUQFrtCfZD7PFs+Y30y2
XgEj692dnXE4vzVY+6O30Li+18KL1PqDx3cNJevAG7WTy14PR1Krl0WUXCfntkRaJBBISVuvz1uE
t8Almj5fS6D86X5AKY4o9F2bZW7EakISXBvjaoUr8kghU86tiPo4MUNhQTsHRZ0vrwFXMYwZKGGL
17uYiOLBRXnzj2XWILMegOMIbi616P6OH+vsDtX8D3nD6uHdNUyX7Wt4qxUM+51nnDnvkqow8z3I
jFW2Wl9QQBIiSXsERCKb7LukmN3BFrd815VM9su2zpes2mqQqrLc+fOo+mOAEi15lMYzRC2NXAyf
PA8ct1pvuvHP7f6/zdcmaM0K1FzA+ovYjXMtH3sxfyMZf/GasMS7R6xoqPgyjxaEdunpehmRkhQB
tXS7otkHnbb1ZyUL///oc8v4tAutldTrKMQUrVn7DZJ/nHOLfJS9m7s4MVgBcxSYz8oAGJduNbTo
d7BVFn2P7VqnEcriOXEBU7+TUvcp+1p46FxL4FR0QNKPSKrJcaJ6tDMvp6jVp4CpWpyVbJdvs3p7
UfmCtpc8bTc9mkczQR7mC5gKxgySnP1k3K+FA6rlGbLlJgmevp9aiuEAW+dtqlsbv31++cP20vIB
OSApW5+8anivT1cY4cdxX4vZda/NY6Mga6ozRCifRTbWYJX9SIOU3PGJgggsGwHK7Mf0HGbpmHEJ
+PjNQAyKqFjwdCIbKPI3KpeqnvFNKwG78nQjX5qQm5mClxMzRckjTUN3giGu7OuoSMOoqehsxO/r
99+HNTkOMDpCoO67iT9UW+r4sr2baAfrBkXa7jd2kSvohPegQKC2ef5GAeqAr4zd4RFTALWHbnRc
R8yhnKSUcQbEOqBoG1JUxPbca2GpfVqrWc6Ny5FvseGRpQI+Lqg4RUicXefsO2zIG7MJdnw3TTeB
z+IBr4/Rcjqk9nsVDbdC0l/V/YMq9xNTr4nsBeQmd7Yy20tUCmrYo/VY+X8kEU4pzZIdDJ0mhB3i
d/ELbxNIhW2Xhm8aLNA+jeDfsuft4wQjpSv7NFsaj9M+aiR5QbdXoPw7SpxtsISdO7/cPvXZfgYD
SJW2SZxjiC3aRJ9PaT5oRGmvfr0DL4SP/aCxXc53t+tCT6HxyMBWj2C317FWr39trl/i5V1xq+Rj
sd9VCzqa2QYGniv6j/idrNozs+76NYnvuJF7jw0/iOp0yzlAbeD+S6ktNbA3mKJZlYZmnMtLHyFv
hOUspzFrt09NN4Q5hxIDEAXMXq4lC7NQm9lBzjZ50a1gpoCz1rogYL8LaBRk9VCDtpGR/Jzog6gm
K0NdksbDr3qjv5roheXg2bEP9BPwbG4eUmLFG3S0h+NR6HdBht3w5ToOA1FDRsR3biGvwkq0d4uS
hK+SNsuaixz+4I0DGnps5i83576uthGHLMZ8K2trNGsXF4Ixh5StUhbFZNy3d1XLkD/szx9TD6uK
ihAhfiUEvkjUzDvtklm+Ou6JUkqUmQXiUgpGULq2NsG+uPKzPmW90V0gKvrKNowvPgonuVbQj1Tt
vLkYHdW+4Mgh2y1lINaBbz7RrwX5+gPl5+3cwAFP6V/2zuDjF3rIG9M/YSOhFmJjc87aFGTh504V
9qd49CBfpWP/YdrXDVPmNiI/RXlZMc3huC6q3Nv1yj1DBHBe85//3u3jjyNvWFOdvmpAtr0yVDZM
B5g9QFx5D22HILnhMOv6Un7/M5OOjjSkyrxV4yyRWeWZgQGpEEsLfi++IAEuXEmL65QcjRMC8avM
1+rBRXygGTrUAc9UsJr5hsluMmBXgpDEelQs3AQzuqIvX9b6vvs9359FUoS1bs+dW+mFnNMZ7TCb
mNpD3wiHR8momRimnKiLESXYDvx0jPG85yZqnSPHJDTYo4edsE32yGVocfIQJ9vycCKmbvKelinH
z2S1lvlLlMpqh6xAgiNbFFPqRhG97+jTO6FYv9mdUm2uaAdyg7CACkyHjHL30dJhOnliCcJUyAYm
Nbx8Yd3neAidoK88Bpvdua1HYd7nfzIAETDp4ymAFy3grVxL7EFmg9VP54AQgXsV0nm7QCZMm2Xc
+Ob0QGm/8ak7tJZ3hp18SQpUqfZlnvIBKCQlGcCO9BKcP3yOSLIJ+NjbJoxyuHd/8PmX/dXBM7Kb
PBtYE8Ugbc+ylbuG/6wLpWRoTQTQ8xlOnGbMfbY1vJL5w6FWajZybKqJSYrzau3Ml4UMUhlG7IY5
92cliG74SWOQQP2bdLUDVUBeCKC78Ir3o2Qsd9clpEhMYqT03cdzcCd5kzKs+uVtJWyc41Ac9dyS
wX4jEI/At113vslG/UPQkf5BN/r4IPb5KkJ/SgxcMqJvfZ97rJbrP5S6+IONYsbzFtxcDNfHugp+
m8ksYLUTqQQKm+kDxlzGGmMuDxYU9L9K0IssWIqwvgWFLsOEjfylMvVQh65rBIZWMY+XS8xzjiXK
cO7RgzyGC3FkbtyETjoIelEjJY2RCrR4v9oh5V2kZxNXuxAqEv8m5Hptb7DEFss1/4iUhVhh68N2
B0DDpP3slH4DsxvaMfba4dU5FomyIR07WH3E8FRA+QTvySf47+8mZdAPtvwL7fD1D5SvMRIXPWYJ
LQQb3R6I3CUVDm/LTj5NnXg7I6evtCVXkVTVUwgS8c3IdqBx+LICSP5XyeG2q0pfHcWhf3qJAt3Y
5IOOYnJpZaDpcZWIO1+raFs9MyfN7zG2U4C3PYzEJz8o6gMM70aFiu5Hg3KL/Sri5qdI2MHhMy9A
H2nJWSWJtgEgvORIDU6eS8qNZek6rogz6x6Tjyu5OveocvK2ljnQ2OaArnAhJ8wL6giNvi561Tsp
18IH7uLN0PJ/bemDEIi6Eg9Lr9b5HBSKX9aVwU3xiOaPDbrhHAb3N7f+4ndUrqsUgch6bk6HDf4e
sXGDf/nEKKOnuGsiiBV7rxUy9b+1uji2eW9qik9cZ5ZD1XLZb1Z3jALeDfRtVN6realU320mCw9R
yTOBitmQKP3VOFHpl4CBQMbK3jRo0hg76keOqPtW5VAHLa2mxBzkz4sxwqgq8j5OSTo1I7F+QdPz
YRqIMNC9AywpVGqNjeuL2pOtH6gqJkZu4Mr+Bnrew2Eq2/cKvfo+QGif+89JDbjZTuHT9MBBtZBE
msWQIHjv4RJVp8sEYHIdP1ZvXVBqFsWMquAbE8y4NCxWGY8N92c8pzfLGTUPoly7N2P3uuvWq3Po
NZwnmSrtuXkFkYP/STidCLHu76MEUFzF6MZKB/2nalfR2Vo1uuMWwFhdODO2FQ4kozRXJYaahD1x
i5l8eMpA7szKtWLjC8LeW6S+Mh9lGQjUcS+UT+Aef+uJtm3VISLreTuWsd2SO8ILMyyRxpVVqkhk
dnMKyiIMkXe+B3xRkCMpl46PS2XxLD1xe0ZvQ50uwe3s0/ld0VpR1Npo9tEvrrDPunT2vhjjlFxi
YeJUGyOl0Tl4K54NsyhrLymrWMM/5U6VY7guIoWGosyhs9QrrAsWLcjUpmx4/ZfBkyG/NdD8AFuh
iXgIfQ+PzJOlQEM+AOqIc/cg3rw8tm2GTu+eHQwT+Osrz0aMwKeNPii6v2LPcP/Picg4X0zRSCm4
ChnZWV6VpqVLunywYtzEZ36k1rZKvdhuvqAKFQ1jg3VWaZHS2iTtFUyO/zBiS3GSDmTOXvWvD0Lx
YYcDA1UgOuri1Ua+FwyRb+3/9PammneidabL4xc2hFDqsWbDFMV1z3jKvsj2oXnYKtLr21Uf6z9s
ay0YVXLR89RSZi7SsmIgLkg702PlRsz/PaTLzAoY13X5ghcCZsqV8u12Hx7VIlQgj+Q2xsy9wTXT
yt6exGR2qQ4SBF2zmVKWJJhoxdn7fB7ZqiqmUYu1QoV+LrD+YN4gOiMgaYyW2QA/SdzYMNs2ymN0
9YVXiUIX7CjnxHE8O/07/WLYCcO8zZyBCn0I0aYE8AdxPYz0hwV1EqEhDjAYoWspz/JYY7VRkaSk
HF8KyeZfyIu/e9b8UGhEsQRboQMJ3SRJjclI4dtTTpxEuImgNb9iPpC11f7132Gp0LTHqDyDUgAX
zrkcdD5Ab1XFoAJ7EIha9fhp2FbDTvHJadYglHjlZhUEO+scvGh9+MV40/SocHgOJnQMBA/TPiKx
8niqH76GsZIRJT+4g/uei6y4K+aL2woUxpRfrmpxHUiKObc8OIJDSETy6IiKPAcdtiYO+nUSZBHH
muCGTdKcf/FlIfTC8eiQhUBbrBszuNj4kHCIbodoChD3HvdBhpm+V27nfN1NKigYlG+MFNPnKGSV
Tpw1mjje3JQtoofKMDA9Xmj3WEpI8UaclME4m4ACdKOcKUmu7OS9DcuI+ZokSnb1f3+/jP+JE0Sb
/fWrFITbOPrUE2UVgF7AlouQeKRUW1R7QE7UkmBfw6lRlwVSsnJwuWvIyhvDwrGKx7RnAO0cxLiL
y+D9WvfTsHfRgsV0IdIoW8Hdwmc9E/EyzHvacIlPOV+x3pERSlr03T4+B836slZfh9uzVUnEXciZ
1JgKmc/mNu8l0q1On1ivMkz5vrs8EPb11y2kAGxMegHJqoCE37hQ0ZJyyGS/AM4jZfP9KV4yCp3x
G9rbr2X2kaRUfAd1to6+RtaeySiTFlTEC87d1DjS6pvabCVCu2OW/RWh9QWWszGKbiEwOqwbJwUI
vxwjdHGQJWHpeisGTkysAEhJxTochO6PXkNV7Z0M9hz0xCpoQA2Y+j67IFHoTfSRqXrSne/P2YrD
u0FK9WZ/vAKjpTrVf1Ml7bcda4P1dXaEFq9aU7eBmJgBw3PPONQnNlzsbEx/GwykwKsnEMYiCu0v
IFmqmFUy8a9JjEY/zFfXvXzfXGsgNMyTCNpuwLUhcYfc1dmjRPWRibugfNkgQhKVA+ghcs2CEV+u
TgqqOAAI967anIq45/SkmtavJnu/NxvZZJUU0P05bTnAGG9O0TQ1ANiEjjhY30s2thaiOTID3dwu
02/+EYe7//qs4mVxE4VmKUdp/qSfi4jsRtxnSspkKmSWh35yVh0PjhVcaYT/B4QsjUNWObADtfCT
rAE4n66Ed8Vs3Ag925KEaiZIKMIflFVNLQQuPlPbYtz7DWMqyuGgccIpcMNe9eiqaFsjGhA+JCwB
fxwRjMQqV8CePrT8sqvuNh/Daeq3dl3ch2A7ySMJu/sRVLNDbkxibvVUc/OGWliRgS6tWyWo2fYa
VKm6S9RFmaFOZjOgTusJTbvYG8N50YL4QqYOslSNKFS5Xyxb22aBMPA7WPxWKOmY1OzxVn4tSZ2g
lb1cDR+PcMGG3/T0raPsZFc/fT5o5kzicfG9xBW5BA7krzXtyFVDCqNMVERVWHtp4y9IygJ3ovQ6
j3tDnQ7t6vxZrQXkdJaqW9MrCFQZu5dwenh1Hdgils338Setgit61ChfPaZKzCvXgdEf/6Tp3MIA
OTo3+grJ0x8ki/EgIyzxuMdkXCbeyuqgJZ1L8+w044X3HXEclY1S/DuxFSFQYTNEEF3PtW0mRHHN
4KK8K5Yha0vfaGStENTb5iQBeOpSvZtDA3edNUiIglwIqwekq2Qf4feugO5QSkVOzCYsJa9zIaCY
B7vd9JLbP+heT0hEGheFjFw/JjO5NqUdp9IV2NYgrmLZWvQmGs4hhdCQRPv1/LPfWajFIb8Ve187
+Megj9ZgfpBCO5dd3ZhHqrGz0dOek/a+0etTt7FG+glsYuQyucjmmO1+VAtbln1nUv+h/C4VeraT
3EoKCqN1AeT0PxuvakRo9DZJM08m+f7MNPEacj/HcW2pf2aq7mIEfj0GSz1GqPPU5KTVGucqbC8l
aLFVPjekKkKqLCc1fydHT+lleguGKyCYOBkLJpYnm8oPd1lovZhCIxRF+HmZIa+TsrDjGna1V6Kr
MmazbXKWBDetBJGiACOgrj9QkPfuLExrHCEIBcXbA2nNXO8TtfHIjF3s6ybJ3Oxzn2jg1iepL4Ry
q67jm9KhndedJKYR2xdJsHTgeVK3fcm+E4M9uQSpk+PJNzqi8HOnNoF2RRqlHNOqjHAD4l9JWwtK
Je1tUCvVgTG+fTQbnVY9YitlXUUZkgXMpva8cHVMfA00TPY48F9cgvFS0Ltu2NzlGeebAogAczeP
Pp3AE8I0sGqOvsEkM2drEkTlZwopUtknafnCmdF1u8PirJpwLrW9BPRnVkoKcL1DplAYiPBqr3ll
7apbnJYlc4Bp5VAdd1S+NrqNg3dUEoL0kL/qwHo+8nj2cm0RBRhYtAclsC16YODuv9f1R0IU2DhQ
akEK8pdOX/vNhilYHnHzWywGD3ydg/XSJcL5uLTo9aVU8/zRi7wUfbzLqP23TLAzMDCW8q2ySxJN
IjZIS3emVe2jAGKCtx+xevCZDUGGvKQGF1UZymnf5UYEYI78SenWp5Y/mwyG5SnBZEqldW+3zjOI
gSy1LfVxbkuu3u5ffx35WLcN8OJPhZvIxQNo4+ngvijjAP93ZknJIuYkETOweqMVWWRRkgiFaxcW
QcfKXM7pkEhgfHzipbx2rrkEx5ZeP7ucRiYkhAPwOzcTzmUOVZRdc7/tGOi//mXd9ZqppOQB58sJ
jbIgnN0h5vO38QO82Vy/+MvFE7FnDJjPj7KsxInVamb9FdWGAp0gAveqvS5hyE8Pm4pbe2E/TGHN
/f1g94Ka99l3NErmSE1+9ObteGMtjFu6usa9lO88a1nU7AbT0v4+a3rnK5Q4pew4f2iRE193ilrK
UhfmxFFgY/ow/SbEzrFIAbB/dNbnBZLPDPiIjzcbOatay6alKmwY7xdb1zEIX2VvzIxfhEeslsYo
Miehs9vKXf94y2u6dZm2dKnHiF8EHEM/iYz94cQUsGw8IkGlAeHaoDBi+cidGMAgooZ4Zh40mMMJ
/LH2AFVdad2lqJLw/vcXdWZGocCYvSbBrknlwONQu4uDbqsW1Cm1BBjka85KN/dktv4nWeb4NSC9
Injq4Zltv4gfokYk4eSMPtpBp7wtfXyKRrY9aKJi0+9SZ75mu0aiN2H50I6xlRNZLyj7FaJX5fZW
2flSSKOoiI4ca29Fyvc8OQBxMkqOYvQene4pMnW69F6HW5Jx3I7r5b8oYj+YFjhdz9mtlkl7PJSq
9BAK5nHCbOFLtNVdj5EBSvTTqoVnz+UsRIWttwb4rgNxB1aOi0mmTRortHvXxYdd6SyFAog9jubN
q2mECSokGoxhzsLx0iCvrq3USGn+Yit6GF1N+GMUByZ8rjaLozOREtQk+nXVb0L0NHtB83UhGU5m
jYiz94OzMHAXs4kLWnqw7XDA8oma8yQnek1SPhTMugkzGYgel3tNNNnfMMlG7AdQGrrYtdg9g6UL
9OPOfgCpdqI/zlFokX1miqAGLoS9ttl7oropaOWqDcP/D2ejqoO6O54vdmHHAQzvVLoRM4IRCl0z
OM4VCcbhar0AE/NK9fUQSracc3OvfdDRDtYhMW2cLwKPcM4t1n5fTMJk0930E8jdho1sCOJZbgOJ
mSSEz06SSPDrjeQug3hPNbMLFlMXXHmpXy+1OL3UXSHDyx5+rnIX5gB6qQldJ6/l05H+fTvW/kNP
6qn1k1xOLFy092zSWcARnx2Cw3Eg2sc2anc9OHDCR1ftoJED9eaOzN1N1HeEdd8BHMqdy+nmpJ4d
0h1QzFCnsySZW81aW/Dx1hPXRib332KPbnbSHd6SeGiO8osV2aLzlcha2VQJQ8Z+l32HNhGGqBNr
lALyyAZ8zrldz2wYcoxGap6avR7uLGwnmaFpNmFO3tfjRSLBd4/ZbVGIwdw+cLbv2HkF+Nl8t2hc
npoQK+tfVeVIh/29Jj4/UQWn7g4qvLaZBlJvxBevO8HqtGQ9zTYHDHe/DEjCMv4XMKSJZW4Kg+xP
r/kyk53DoMCdzMAdIMiFT5Z8rWlJlavQjY5UIz6J2WtnNWt9Ad68JKdNo05PmV6IfOJTZRLWqAKY
yPgnxmU4RuYMEcXyQ9wk4UHZLduza2NE1sXkQXBfKYSJyHja2795MygOinjVkUnZjUBxV/qw+p9C
wfw6t26mNSuRAx+jJ8GAfx6D6f3tDVwLBI+A/aoTi7YODg==
`protect end_protected
