`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RjBOnpqHtHSn7Th98eHEXvWyBHe3T/gX1ti9+oK+DEEpXjYJihGx5qABFhKaZ7HnG7jWsuBRgFTw
VE0K5T9mAw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AD8tLEblaOjB+faGHLQIkzbrG4aM6nCBT8dcD81Iun3SQOUijB8ABDIg5lEYH5K3EeksCSGHki8g
OvxbLFTgjliJBLxLsx+ia51eHHbkDhVrKKZyRVjuRNVWUvpPqSQue0dt1m+8vXZ8EbDTFu57FQES
ftptMOmvCz4P45+upgw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Dd31zkgUgmtbPfI+NIw7WlVAEr8tSKWNShbB1sHb/DVoeVc7e1sPES4YIchOZKIfybkZs4GbQZzu
7p0DR6LJViMcpdkP8L6fqfNzF1OhTLtyiyODjmJKVbEn9K3WIpfx3cKfr6NLVyyNtOZfkBdGi5Ju
yPztYIemvy4+HBXWlBIbtGcnfXdNFt6Od4zR7R7/HusvUvKc/AGqJmz7S3809B2hCVf4LcEqkDzC
l8O/4DarStZq7ROZLBUD+boey+5aS2clMyo0UHdNPvD6k+zdaj8GrnfawU2PU/hDlhDX4CeV6VAR
YUnkfC0yC72QCfwlKJ4gUttkmO+HsgYJkC+aOg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QhWl9RMPJdD/ZzRR8EMwTgTNuPOKRQrQFdbwGVDvZKtpMwRqT9R3LfVWtbQcz8WGEhjsrZdTQ2Tt
VXYvZIIO7sMT53lhA3efDgr1bk94sKVKucYzrMdSlvkj44xuzeTUMsmVRrIVvGGtMytti17Vm1/W
vosV75seV2FQGB2C4rv4he7Cogzs2UePX7lT3jCmXP0VH7iWZUx7ew5GrP2Lte6VI+nAr6bYcgvE
vgA3qG2GsLNZpxxVVGWNesA3GqSc+PIUB2xPr00h4vrrgYxO428jrUtnAR5wwUZw9W152bGVgIX8
xZau1x+uZ3yzQTazm9yu6t4ME2PBCwXVz17jDw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jpkTKe1I/bpe85OESn4XWlnPzxPg7qI9WIaK5XaiGGBGixYLwRzLlNkUzErN03b7oqURMr88K5M4
jNn2+jzz9HmzWdP0ZGKTlhrW6Sdko4T714+/bxB2IR+v5vpPzrpnI50QFbCjIFmAS+RzojYfVaSs
9AwUQ1qyecUtyzkjygo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FnnZEWGd+W7GPfbxXNmL25gL5GeM4EahuG6OQnjnqdruSkYjP2R/neKgChYgKz0laVTQyyADbUGE
HLaB3cP6Mshm6TnsnznSYK3MYY8w1lwyPLH2P3S29O1EOQLfDNE4m3G3ihbblMd78y/8SmJiycPk
go89UvGCQbKY9DEXc1lfc/kIKXgMkB/CNdD4PkOcSDb4YH1FlP8KteLdVDv12i1cLvqCVQYiZIvr
bPu0MglEawi5DZttyhu7zb5dLJqPtl5YpEeYPpnAKqKQ0+SJhzfzjc9wrtkT7vf0NhK8OwYDgbp7
wX8Dma61ADq291MJDKSyxgY2OiH7zkhHt9mvdA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k9ONE6V8cDPlTUs5hhzMJIw+J7u2toMV3xjrlyeyXlJat41nqtoIXMfKe4BvqchMuefafW9o2L9r
11s6BZl20Y69RcOU0WetH72qfd7/7Kpp+ikXD+VrFWxzhaZufypkPXMtQGr98S0nR5j7y1TFJIJd
qDRH1OuRhVjJcgd9KVnrtLm9mT/oJOOeiqPMHaqf6aQFna+ZSigYPN/QMMnTMfSsdJQLmLWo6Z4/
lAS0efB4bdfMEzg55uYjJstVlH6jQr/CRM+9L6IkMoFxPYHNWqS7LsPs/zw78SU/JnA3/cVvx7Wy
RzBFiRvPRFB7x6tSNas53jhf6lVanpPxpin40A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NJ3AewbGy/1b3Q7grl6l3g8U/DqAzeMvF0M/rx3LiqYv/mBQyl3As83UPy99ReUtnyfJP3CLmF9r
4i+XbKr4we6uYQcjbnhylwEw56pFm7SGXVTq5roiDHSotdKqcr33xTDX+9/auKrJUcx1Lf5rScgw
m0oxolc2QVL1yT4tMLK/R4C/mdARmD1Jhf7hKfUOIKi/xNXzXcqfBPU3jQ9AuZW8aTM0nILtH3XA
ZHBcPwZv41mguaikMmdwlA0v5KQ4jHbnOftBLuEpvG4KDiFFgCVN0rxTp3ObmKYNi0n/sIdyXwyu
xJkurQJKLU+73OaQuBjToZKkK8Hi7opi24E4eA==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J9x89Uvo6pGaqNI/JxQkXmn17BeLNJdHi40iwXG4XmigXrbTK8r0txxMjDZPf7lGcor6U/li1IgB
zqsF3jG03OqOjPVxJz3ymVNO2uLbm6Xefy/o5XhmwVZIwmxxNRtZfSeFXJDcLqJ1FEOUpKjWZc9w
u1v+F+g4pKLsoQOSnFRGnaRfLErIqY+NuyhvRJXNncy5oAd3mY1c66jcpNLqMMjIFG4OXxB+NeYi
XGI6+jt4apOfng5+RGiJVzA88WHZIlLzqgXaKg2TpgBxodNUl7nCUIADd8EgIGdiLaX3GC+IKIB2
1UO+CctB6E21VKAqU74VG0lD/p93HxBKnKjD1g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 261328)
`protect data_block
jzPEMC1p2P6eMSuRFSavesO+G+c4aRpSQ4mybmcYBQqweYgtwNt/k2WKAh7Yoc6zVjiatzRb4k6F
ouWSgTUqf0yCDmST3r81BpaxoX4uA62F3d7gS9dgeBRIgGue/vBb02j1oO/VqmsH11so0aFmyyUH
V6CZAKfFlFg73EF8sd8DyMcgpZFSm4da/qIpb+vIy1EYat73+Ux44p+IvI1npj9kGQgf2EfKUfYa
w393vMWjDa87sDJl5ptd2pdKyhC2ZiQk/ltV05scDp6z1cbeRHGkoCjGgPSMKW8wcwL13Ho91bli
QDZoHfVbBV+ZTssQXjvzP0tHiEZs+t3VCkXdcFZYmEwBmYZU2E0Z9MLNekjUd0EHG4wiB3mGcxer
AUaDqRkGtgMe8fhKEmtw/RCLHnWFBkZsoS9jwvcfr+PgseKPconRbw+eKVei7WMvC3d5AYH5Mqrs
FPMEF+2WYyEYxTMl5srwi0KBxEAbDN/0VjlRPL9xP+n6XiimVeq1N0LK3jAoeKAmfy5EcpxP5Tk/
gdv+25nPPSZ7oUq0L4dbNsNayAhZgW45ddSqhPZugS+UYPLinJMkt4KqAdjzgzwbA4ZiAVeBku37
Qn74vUXN3Sa8BIMydGFCZLQ16OeVlgUtL5HI1oSEobjcVsUXQd6ZOP/3OyTJLJ6EolWxwkFa2TQ4
QZHyrK/4GA79uS/i3oP8jqkXWK1lXTZMmIt8Puvqgs2Vnax4BdF2q/wYDsYG0TsEC194MmVwDk95
o5OUELOIKo2hMahx/rnYvZhpVB5XQo4mvJ6Kcq+pF+3J639GHvWq5utg8+EMKDtlKjzCgG+ccIZ+
VH/R7WKAjrW6cxUmU4OV7gQzUcO5ieMX9meFMcLhQ+b2Mv92dwaxu89PwKuDRmYh1ZWuaLnytBdw
eyEhZR5zTSdqgV1TLy4WB/abcul4SKJCtgEF65zAtlPRVCHBsYkbbAfvUgiTWaTkI/fCxnRk0kF+
C8f95hLMHn57MsT/sVU8d4sYyHg3M05qLZiSjnNXwYEbIYpAdIjl2kJOIeWNGUYyucBRdV5kpdsM
S1JPKsmJFgcH3BIaRnonLXV2Z9tDo0nd2GsLRpbyZ3PCbhb1Wrc6q2mOlaPR6Gradts6U6B6zMCo
6cXcoxIGezvXd3lL67COXxmUzNdFkadLSv1ngX0zkb0SB4ZsYg813G8T2SASftCQCcpa9szq/Qij
N//LpUX4w0HtlBCK8YEg+4f+c/2x8p7PUzTXo7ur8KaqKgiA93L7p10m3YKQ/vRdbtcGrEHf1eia
ct4RZhfjNJ8/JOxGg0hjYd7Y7oxeVEqg2TFI12rytIu6D9dKdsUmo96MQRQqYWcV6vTjyOgom1B6
AVf3nhdd3pwcxhrqcn/FDZstktSe3KjO/lHA4NuicecEic1ON5m7BAZy5Q6F2PPfBtS2rEEGX34T
6ewrXj25tBFr4igIvCCBQ+uQ/orj6l/hXVGaKMw4IKIzhPDeqwPMomWwF/f62LSWP8LeWvcdAwQ8
wlNc5IyGCiXL29Gbe+j/mxfFpzS5WHzEJKgXw/bLyBYSfHzpxnzw+V88DriqZWOwSxs9DVUuq5+Q
fkW0p3q3pwkJMa9T/XIObssU06Eokt4nRIRRvcuwAe0+KkAo8zCZX30d7BxFciUQmQ5fUaSJY0kq
AnPNzmPGVdXAlioms4vJLBghfz49r+/3OmHuYCBIqWq4uyGWF9uCSacYRCIxLHrqoeGbXwkivyDA
i3E1ZYO5etA29W4Ch2NxqhlkvG/GHeZu1YPX0lV/SXzti2byTGDHV9ehYSlt5zsOPpoPu2uRuKrR
kCPVXH9cVdhAlScC617zfTLtZ+5a5nAo1j5SGBqnSidVJtpg2JSH+AqAPObsXvVfTmWMi25DkStq
TAhGkWrWer/Ea0V+YDLuseUH0n1BIysc49iipg8FRbRlkYq/pH6ap6aZlmgr6g13o0e6vN4L43iu
dWIEy1xOTD0X6L6fKZm0T387H1INmaZVg6npQHnI5SFImFP6YiVWdtCQudiF52L6JT2blUvU0uZB
+AtVyT0p48/80AhlnJdUZxRXUE2l6WAahFQw7lHft9gbA3/uxa35jiaCp/v/h6duuBicdDxdJtU/
9bYUGWapI/ABA2UIHgsiR8ZdAugBouot35lV3ZYWwPqbkdEAv1qOzJUf3uj9+mRLGk9A8r9G4uZs
6tqzBNqxRXHQvnC+6jA5gtEGGQAQ+s0N7A360NQ8gr1Aoy98hyK7+1bVCwNeHG699A6hY1URKVW+
S3ZjGLR7CWKHdiOxDhWLPlDGjTmDBktvzCq8mr0J+xRHML3BV9p5n/Oy9C+HcWZ9kIaRY4/q8Sk+
u26dNmQGPUc9/LsKmZtn3gPbmZDz4Wd+lexvasgZQG/EVYz4oGXXrvEjj24Y5oG9SYjf1jc6iaD5
skqwR6MTEAmdBsRAXW2AcHdGZSit9oxg/WIfWelYzAHjnI0Xcs6sQ3AEJ+Ob1hrEi2P4viWPP22X
0TkIcX1IyWlVPeIUuiqO1ug2LbEHNAZFvHn4xxABtKvx5NhK7dp1//bfeIkUDseHA0gQvQ7FMgPM
JMPPDWXie2+B+v2wdukZaYbA/rAhnpE8QPxFjsVPlnvMX412Q+7AkSpsbF2JVt6aBymcbjnfjYBS
9QSR8tsJOGaXlOhK3WrXJ9Ot3BGu1cqPiMvexYTMD24wIitjp9CwMfa1QFQkAfgDcDW1li/SsY9H
RlFTKbxx+VI0813IwxGuzbbTm0nnrWBkad0w8uS1RLyBVTZW6QZAsrd0cfq4SCjX7j39balaD0MI
CCIw0Xr7QWIfhhgAwNQtTNpHWY4ovj0U7UaAJX1FvaeDqYwTA/uinSQ/3lxogsGpt7MvXGYVhUO2
c1mxzOv/+D7BV9z7y6PRhCvX+4OzMlAlpWC5oCNgw0VxOH9NPi+y4pK9zTsJG5ENmZWRaJ2AKZgI
uyTcrSJAkmjFaavER9l4FmN7njmHCZO0wDCEWHw+/OoEDi4ZGacT0sAd6ChEgzscW6e/r8QXdTM/
q6K+AwfWz87TNvEsG01hy+gT31uSSD9aWwDoMfhwLM8VwXjNYnH7e1241CN4dt1XWaeCfWZbYF2i
zzwv0+5D0gpANFlqd3cBC1KtfKt5r7119bbS9DzfWT3HNQL7xQO8RFp7XEJxMynwu+zYoYguSLdL
/QkEajHrah1DLwaW+unF6E1bhV5bNOaivEKRFc8Lr9/xvsri2Kee7VYtz5UG8meouYlZmqIKpWpu
hUGkg/2Y4UERVrXDLF/ZUGQ8ebzCgSwVni0EtcaYnd5dyeO9AaXMCLaVaQyG4s9633zTQ9s07xPv
vxxtlGAggg5uvWXne5fAKhxCOEAf9lyh535R2MWhU7qdJ+1PGw/BT2k78crSOHe8rS2tJ4UySUjg
BeQwsOUZArC8WwcuI/o+pXNqfGBqlUqYTCtXjCjVNSGdckaFmDRMM/MuEkU/YnxHPkXdd/qmojPK
8tzZPMG65oJ5w8+yNa7hPeEgdPGt7xHMCqmVbdtjCMbLLYJocofbSM3RGUF/32umK8WlRcd5eovx
FJeMlUGDgEjjeFMWQL3sBz+d0cDrBLmbcNPMEMWzuZXsrWJg5A/PjUMDcw1MPii3G6lDjsjaLUXY
wtVuzkFIpLJPz7Qd915Zl+zOdCKFpFT8CSa7rbC+hYLwPpbT9RhrKxDbv+fsNHTTuNpeHISpejVE
FBQ0zql2WBi674ycFlg6AXDmE6ovJzG4kfD92Q6djJWS1MeQHoJz6DR0YLd9bH/ckLr6QvcXJiEC
YGkypgHK3ixQXOHCPRPui4ogS6Y2egNS6a1E2OKs1ofOeqFfeu92oTptQ6O4rCask22ok/lPwOti
/RokWhi9SN/ZcuHq+i5JofbkiCXqltyz7PFEzmTsYLJWAfQhu1mzXh6uh8i2kUvUeagdYdb8BCXe
V/dCpvkTbMsWlq/eBUb+D4f6OL4cRk7TfsXG8brvuYfkpTu5AxcbJGVCIhUpwqIbOum5zYO/HtCE
n3OtUlMryDAy8IKJyWoUawUWeuU5YdCwtuZjcicLG46HNLJDf9J6dP3GWXc0tXwnonpcRfHXALZl
1GXHKauCPeDJsZr0Q4/zRaLGbwnDSCZGFX2oeC68e8KS07Md/QiUJ3cP8vixsRbNUMeuCogsTrXz
ONtAfwoEviKKsuIi/KBF0aNGIOOv/fQu9Gkt3BHD0lfnFWJ6NhApXEBaI3rABXixWii/31XaSEhh
6PKOSWtj3GXrIi8ufcCUWaot/EJ9pk3ODcF2dyxk4MuigERPJmAlegHLZuopeUkFgEz1bADsUJjP
8H3LdE//BjsYtLIZoWqVcEBYqfJH264++l78tAkNPy7Mp32OErByNW+gBATP3H04XWI48MhV+UBI
DwHAvuKN/LEIuhpN//cnPg9A3YfW69HD1nmrJ/StMqzZQ/Zzzuoj7YQ70qguID64IMmiVH4zGFap
lONuCXUqV7eyjIDSpCgbLoVpHiwCb5DrHV9QUnC3CcPmakj5Q8XbskObG475qAYJ33dpQTvU6YW2
z3h7wbJF+AHacU5QHop9e9/hk6wDXSip2UTWSqh/T9++YdqQPTYafDpEIWA88nWPtyTEYV/59/PK
+KA4ebOs+brNLOiLn7w5Y4vRkRAo5EfIQkUWCdYVxRM1hY96enGfY86OWxfZKnVez/ZShvtX5hDR
xvljt81Stwh5KkvbmjNpRwa20yNcCD55ExWXdr9ns7+48smk6S0HhdSvMAIPKNcCrX0Gvi6zd+2Y
qI0gzTRiBaASuvy9JIeXuW4A8rNunZxq+rCWsuQn56Lx+1aq3bD2B3Mx/jykypGjy3gMx/h1y5jx
Ti/O7qhCJ0bvB7YvDphJe1lW2L207iG4uNpHXIjmJn0gbSeucnjNYgDR5t+IG5Gpb9nLQTshsgmc
ICqcaj+eevPjJ4n1xfr5Q+dxde3UAEXsMbqjBRBVdoOmkKGjw0K28Uj5pvXApa46hszTnxBLzEOb
esHN39LdBQAlpMY+37TdhHznvyf56PvOIAPL7IwE0Do3ffkT6geXclaJr4Ns8ta9a7j9NNKcjsbl
xwOGOmsoYZ8vIxjfdgFIEeslGvZ/aAZydKiOYn0viieefpGqBV5liR3TPYPMM2/fDr9AqfuHg4s6
x7Zv+EW96fiRKCJmYQtEJUsZdqSOzOIssRWJucaPpaFSZIFhYm6ESkukKgKahKCwpraGF3gMlBl6
ZEakg5Ek5hP1SNbt+GR0He+RPfhZPKOyQi9wptJuTH69yyakvRcr81ylOLIu3pLTmVtsVnNiQ5rE
3vKicweOuQB08vP3pqjY7JEr4CxUJn0D1jbEt7SsOWns8l1FRrfj/0C6f9spryUXtfMsrxjnWSjk
7Te6WWdDdxBPfjoA8kiPZMqg3rmwW1rr+6FWI+p9oPs3iZva1X5Cq5yhmyQu1iGvBscjdyUo/mhS
Qs/4kQ+2j3nZhUgvUg+cMrzAks9oWck+5eJffBPvHBF4zRe7RmqV9Apid8YaVon6NLWIeopuC91x
QPzU3Q05z/TjRr0Cc7e7wTAB920LOE1j94t4cNVwck/1/DsB8R6Bibq8QcYsOGoqdViYtjxYlgKC
erHFIK1v8XNY9jz63hQC9LRUWYMPeH3Wl/DLuCc8j0PjqZFXXI1WsSWfLdWhOCmg7JAOh3O26O/Y
y2OU86TkXn7LU2DPZCBxXwYolvgDT4+JkV/ua1lvPGYoWPAv7TthEjnRYHM4p2yORXqM6yZ+79Jc
641ScpwsvTgq0LTVuxNMtT0NCG4ZvfDV3kDiXh/V40XpD94CFvlr5++Dq2coIc/ypx8GMW4at0Um
hEXcELzzOOvZtzmgLRneRbpNmI2LhsR7dNebKV7C1mWztZsNVcktGWkG6SnvZlRr8ihs5yqim+KQ
6mY9kOiNbYb/K0r0S9FZ406+YHAZZNitpfDMeptkfhRxlkyDVb2K/wpx1wA/TiBnBK/pnxlFkYwY
TC9FGUwSajpYZm+SzRl+MaYOFAfG8iXuecIsTv4CwxjXI7gbx6e2FDKFFFjZnkDKMhvyTt5UjGUn
je1uN9rv2BubShvfyywYIy47zlV/nWipOhhSPR2VTBAh5yhDzcQ4GXWKr8QF+kF1DSeIQ7lSbVz7
iz9heYmBi9sYbP8n8Lr1JoIOn0unCq1KU+mm5XLDB87VQxQjSJUyUQ45/1OSvRWR7NacVdEFogQ2
epqESlUk4Yo8YQWnA6HFAdx4KwxLuKpMstUA0YfkJV/lBSJglHK2EL2pqnrI9LKWMUmHvjtZ+qeI
FUkGkw1zna4WJ0UJlVUSXyN79TL2yGmS0DPMO30Lx8Gse9zzTHkb/5rUEtYDK/x+n1efTjeFkgJy
QIC+fbWdHMuPQuUnpe8apKAOIdOhWbp1K72ZeYV4uUJazItmkOQ9HfYvcfZIDIMqXpxzJcqnA/nJ
+PsIIjV47XDQyO1J40PUa/1qvqoIZoLRrQ9SJhVeI29pk496HM9cg2IIYaUgCkqJj4NxbMSlKfAo
/2J8GHQyjsCWlCPTKfHNNMdroOTD6LyrjJmG0zzIWzBAb2/w0y/8PIizDPkkNGlv12O+cJrILt3P
Ft/7VjifZTbKqAwPmLf2vUvyikZj74diWZL7ml7TddxHSRWd5cPyU9pNwHhlVB9S69IxRB7VbMAH
oEAGCReUN5NTKZMSf3ABiHUhqCKvlbivq2X50msTc3WlzzeYc5Vi14LFY2MV9fULnw59wHfJMd1m
+hdTv7qRMqSj2k6GW7FAduJM6JILXGukx7F2RKdc0rvT6sO5EeoI3sZqOUnb/zkp/Xj8jnnERo0s
N4uYd+DMSl19v15/me9/l7zuDyNYD4tMn5oOMdnUaS78cyFgV8I9pe9NNixdmhZ5z1FJujQeqVXj
bPxVAMSz3/NzdeMxusidlv1BATobsWuRJ6ZJqXrRvIiK49qMtZtMkE4jBErHAvsvudQmlEB1DZjZ
d1+ERNcx8F6z2D4ovec6YG0Jp0LO1VbUJ/Hs5BVDexDg2mOVMLGUNeTaFrjMJkYj4p9tTIJBXKEQ
wlNOYCO/xrGdXdjQxaV/jbQFZSWhM41odCN2+nyIfhwJg6gy5ppHuiOztl8uFtZUxoBQdEpz0KDc
fI2wHSL4h35Xt+pHMhJf28TuPumDn64TML0zWfL/15skow+BUmfzcuiDvA+H4klFFx2FICkI4iNE
bT/U6R9ivXHLJI9VJToZ1s0MuaGpUW8C63L4hy9npQZxHvPvX1g7GDVgXcBI6PY3i+T42bbGJFqN
4HZ7NOYYGtLVE8zvYn6nPkFY8t6u1xumkrz8bD2QaQPnfQhFmNRjsEh6Hwz9f+vnDz6jBfR8JGxK
/e4eu+EXkXBPepalRLeKV27ifV3A+P9niSpKD1MAfYJpGEm0Oy7Srw66VuJ8bMmD8K5Qu+o8Mvfl
XOEftkn1LSkifEixiLNJiKzfd99VgwwibAYZ2yfDxUlrqmcRie5yvBYA4rnRriT6DaMLzBkaR0aj
I50mCZp1eZNjNDzNXrBBf+cJbk5tgksEYTGdDvyfRMuhj48qgNOXaEGJIdhEOmYqfYneoAbACFiF
VQlJwpz/g0cjnSWFhHOLxyHTPo31xhxTPL5csyyI56D5KWQetvTqO71Xad1QNjqICxU9PKl5NtpV
s+WjfGLouTqbj7fvGZa46wAUMR1j3I9MMbJunB752Pan2hoVRqw+mlhQhuuw2Ml1YL7nY00Yrax4
uizOTz6rZCA2Zv6tbk95jDLES89IEh6FXeYyyaiFBQF6JqyJ3SWjGyux7RCyJ7gRLvq9y+zF1V3Z
Qk3/zQHS0v/X904g2Ckx14vYJIwFph2QyywfkieSdpv9Vcp0wdNaEDscEuu0FlTHiEQuq7bCnlBX
jqKzkny6ypFOYUPXKz+FTip59pNKAk1WQ++pDQChOsn6R8fqG8hZyGlRz7RHTharNdMylyfxUHv2
QzGBOUTo2Dt5/c5Vr4S0m+yaG+teB9EFHmzV5RHm02JRnbYV6tXRNs13e9O5JO6KxeF1dqm1KHOU
MvGIYWbSPuztgNW5LwXUIbUYF+fDBWM3CN/f4ixWGI3ycKjS0CUEDYxjt1HnSHB/ULg0wpM+rDo6
Zrbkg8jOw8PWTz78BB1Nx6SonvlhnE6xxPpmF9jQygVHG8ruyfZfA+Pb00O/VOr8yV3UuC5BHEzh
vlQGXjikZfcEnxfk+vVrbfEPYQgScQMOEV3f3fF7L6VrMuPmezHxDkkXqTd4tL2Db89nsNdYFzKA
ISUJVrRPIGfIp5OYhaS2N54JS5W1XoaMpryYAoqvt7FTksKpHBpmeJIEbN7nplW/8hUsPqFgpDlE
vqO8OJcwWIW2vAp+VojpTD/Xwe8UpS8Gdqe4keo9pWtoaTr5jqxrRm/DZmYMLPSz6CdAuIs9Ta6G
f92lFStme07lo4ZHqusatroqnuBTD/qGT50s5MmW+fgRuaTbaiKRrsE8KaZWBB8BAYvRMzkdgUMN
Zp6sGJ32qDHo2mEYRD94wc76zl5GCsMyk8eUMWIgCQl+IihfuT/4jv7qBsX8swxL1WD8mQumlakz
B0l2sZmORI/PqGYmBAQZdS3O2hZinIVrUiZgBehLi5RB2Te3xaCcuHtH6XK9S5xXo0wpirl8VDR/
8Pw7CAIt+SrDfs4/ObA/WwsVTeetq+yyJBGOKL4xxCf3AnQA2EZDiWZYXL5oz2YpZJ8ZXzd58wdn
bLGgJonvl2vCa0g5Chh4K8nsg7kNqI4Jrs+DTn01XNIrefpJFxYHk7qRZ8E7OTcxxP9zshsnwqGT
pmeT0SoTQ3MSvfr3uPWk6RuCcbQNmMWFi1y8OVZ62vHFlVeSfLBZvAhh9/LeipEEH/OwxDFCox3m
Lqf7PLOVG3GyAioa1mdez3GZoixtgruIVY1cDkQiho+daSbSy93J5X9vAfdkwZBGwZzyJIpc/GU8
Rvy4MXIeBAmLKeh0/Tq4EYzzXZl4SUWAXQmQSc1rAmzQQ4RrElefd8VZAd05Q8mgj4zMWqBSdJdW
OrgGlJA77Mpa9WauAGzD2pkAGO2b0cs2GCgokZvxHf2UZ8JY0Ytvw3YvJDMNtQ4E15p/seOLOzCc
klXprmhbNkL8d5vxg3c3hjBP7+WfZqeB0bPv9ATjUPpbfR8IyRkZ/YKx473VsjqbBPFC6VBOIDaT
E2QFt0wEUS7LtcTUuLYnA6NP+mDvS6wEwCdqfnfXM91l3HAjDnMxUMJliij2beymV9npz+TOdkY1
V3ZOg9grRPrdwrjCc7cs6Rukw1LZzvj1+fW8gXgksNnNzCrIkyfN+hPJob/qlKrld0jslFyz/jBC
wvfMVp12WbaYjoFs6UwIIXsW1bS1ytpZTyDCJYvbDvKP+3oCrO65ufVxGDhfXK75Qlt1F9o7m5pe
qnlOxsGE91DiepRAYW8sOipxYlTOA6iTFQmicO4oxOIltiW9AxHpoW3zydoP9L7cFs2qStIRiPcR
uZ1rO+L2xxLIBSR5xokPozkIJsN6TUT2wHQREv6HNzv8+4JMCaZldF92YEQ3jmKSMZk6MmuBd8kk
BRek2a1xmSImS7N20KPkgEQWnI7fDTubDgE/GQaSKGctWqHO89kxKACYZoR6wOjbM2QgFkA7FP76
RvAdC4ZTCOtay9FzkEdIyt8j7V0pcx3CC8R3FC7RUC03BQ4Hwur42NrL4oV3qtmpG1/5Mu3IdBvS
RlPBxhwuIEwBO+AQEpbG6KxhDVQWdxC8a6KoE6uaEKu5P4mD5D1iWdlGdhAmp65ws5THgPic1NdC
BWDQWIi6I6MUqSVwkcQxbUkO2f06qssNM2BzYMu+WxVMC9Jfzk+0DsZfTfANSmgL/XsvITQF6e7S
MkiSNlKffiKYSh3weEtBbQFK/Yk98ovyGE+CqSSMtUF/sSlA/Hq3ptVGaerfB0+tbBuYRztVh+ul
f+SlEm6wr3AhRDYGhN/X83+6yBc4eX+/JVCuQ3wMyRItg5N57l/LGhS5Y8G+vAk+uf6JbC+hVjby
vzYXmLu0JaVFCfNubrq8Knwh/9J0Im6yHzM/kXtpom9iCK7XhCFBPvSkBnR4cks9mLq5IgYUpoXM
jW2x/QgUn1dpCZoPDSBQcQYdnjSJiJvkidccjdeUW11yKuAcYqAGQAl4FXGOaXMk3w/SqxIgOCyX
UWBEfGOyp7sJKNf+ZUudzuhoZ4STs8dZOtUIYRpWoKSaf+4YUMjPh1kVr3Ra54bb/8LUKwsmiEgf
D7Q1YbqaNNbJQ9hmHASTb24Z9Cg6vcxTRQ6QecOX57FxLSpGxJf4Vqosgtauh0bKTa0JMvuFgQRe
0g91C961kH8c6INfV1UoZ3RMjHHoX1WQxKDZxVCVl3sB/kKE6SIqpesom8KoNPvnnOx0ML/9lJJZ
6UFthkR3jPjkFd+SF2n0v07PPatmkAINbSTs3ENgkSqPEIfKT0V6nk2OBUlE4CagPerbs1dZhPNP
CsYRrYaBz35FVWodug3fWtYgFNi8wBJJ2N55n1bXvAREBYwoYzSHnDFzDZeTPwG+PfsLLKr4/0aO
tzrW/yYt+5iv+99DSXkdINGmS4JlJU6CvM4HCLybSuqTOal1UCPg3qiI8UypyAg1XKJhXvL4qL+G
AWoPAEOAJ+D7s3hLyYFvWdFkFEfn5xjSi050vwfdeHydVN+2thx2BjVnk5FbeAtqprZvV9H1aFpj
J33GvGyJCWKmvbGQGJ4nB1eYMA140GPH0mMT74QZlqUbQmNlsajEEKb1xmKmE45DE376OPcw79k3
Kk+pgSZZuXFd8oOA37/lvth/xzJTkXfU7v+8QDJybFGDHfoNljUQgwqOhUJFXw1f4X4e7W0eym5L
IrAvvqOYIcezVBTPSR3BPpZl/EAUA2YgP+CDIkBx9mRz++nAM5W/Crc7gb6zs24V92WsP5bnI3mf
Jizo7Wl+HTsjnCYrnrMedONeUfEvTuIaYZET+dUc082VrdIKO8mCz+3G6g5GiB4ECn/xnjgJFwkc
yNsN6ChsijsEtF0PcIDDrcaGYpNJrcXYJN4EDhEkOXixHVsApkBlpU9drhLfXcF2UsoBlmOTaFG9
nLyCDEY5Gjy85fbP0bKj5XbmYuKF1iruaMWhLPIuZO1sxo5YugidXs5JwTbePMmj9VNcXzmKsW1Y
FvGSVk3NWNa7xbP2O49Ep3EvQ20/gVg/ZFxLaPdGbxxZ1WdZkAFj/Ffjk3oBGuZ4zAVyXXJ1dYFb
p4fm0yr51hHb/FifTb+p75Z1cr1an8iPRM8/5xBsdA/5aCstNQc3SSgIC9gAsKejuyquA4PRR4P1
uh+cKKgOgiDg8ZPdRVALDvj0UXKNCcp9d9cDgWw00Ovhe8x/nIsb5li7GiKj/pFEaw2ebFi3RMsx
CCToVZLGHqos6OuiN0iCaopNULwGStmIlpmczksS/nrBWmD2Q9NSrFldayOuIodDxIga+5DyhZkB
wo/GWnKlj3O2llwuM+mQ1v1+G7/5S4IHb5dj3mwn58ctaQ0wEMOacAl8sXxziJhilKYp7SGKiJEu
T8YCyNKsHHma+kF+gluDs44PItagqRSLJCsPLyCl70CgRXiuaBme2BN2I1huA32wganliUiw62zf
NS/3p8VXtH5D+W9Cumm+u5TjT9XNcQaxRCK/23+MvHw6osYkltdrMYSnM1V1bgB+qDYSWq5UIQrU
d+lEGtq/nHBnZrvJn0qvcSoM6cSrEDB5zf+wIHfgBF6BNxZgeGJz2yhbzdyNORAlcSMr4Y5+zwRs
K8/HvA9y0WCkmf5HSWMWzZGGYrFjmnk85Lv4ZEv3uz8RgZe9/zKwoAo1tFCFr2fdEdTwaZ08Ujq1
tueu6hW32FnlLGdGA7skWLSh4r5IwP12RD/Kuz18zt/fhxFiZIOP4HOHZ0dOKWbI0/trvpjsfnRL
P/DBqlJbf4ZxXsaMQCVTelKcZkGeM5lUm7xVTbIC2Qk2yiImGZCHa0fo7KUSD6pRcWBFTFOv/CuB
UlUNl1L3Z6raTrH8owYAf1mJd9ey3hIxn8rWyYbjFDrpc4nfRY5A812OAUSq1wPntXJIVoIBYwse
HVaqYSBmga8rh3dCTXDcHJzqtL8paZiDpDu+0bK0ciCkS7//SMCE0jPUzqS7iAA2xEdPXADFL5ws
LkX9p/GqCtjaljvBW55fkm33gxuAkjxaCHy4sSaPbvDWycVQSMtGdSJpUOu226X1Dqf6H4phqm70
eiUYb1jB33i2bmU/wu+dAAWOB4BntpQ4Ts2pgmJyDs0On5MVONo3shdgqr2iqLfCLoZ2gyyAXurD
lU4SkA2Roj0R2pKEIY1Z0ZwYw3IEslvB6+PpjSbo7YAY33FHcPdIFJ/9Z7aNaHpXvdasdN/UlIL6
zQ3XJQoX+lJb0QPIo8unK24Z33/V9/hQudsdGjx35bmAwDgCMqRHT0kGjqWGAI1fzmA59t/qN/Xa
/r7V6frTBF3yB3mmgvamRIJSrGP92/ZZFQ6PCKtqK8uVjZRCF2iPFw3QC5fXDXkDiVHI/WWqiN0d
y4Tqcb3ESohMgusVIpZPanVPO8VLXf/9Za6zBbGDDFFMhJVBTKIMBxE3ifXnVeHZlpLvR6SDdZWx
TdO5+r+xIN7Ylgg/9VheVYzNQBnurT22B3TEkAGHNIV/O6Nyuc+lnZ7PQtKrIXTBeR9m36ch3xya
7voGCtpDdC5+AEB0XJw6MeuAJr/TllJlH+yGzCSvrxL8zitGBgzpjKDAMjWtcEQy+iB0IjqD4qsc
4jSlz0uLzXPFdt0WpfUbXrq74Xukmxpg1UtYyN0IZWv/FoEFEsAh827Dx8BWEywRKxZwsDdPiza/
T5lzGLYF5p3QgZuCb5OhZ9w0elfIlc3xrqqXuPsqfMdZrwuDkBu7UdijdAbgmD6qGhClNct5K+bd
GF7qdHhUH0Qn4NidrjqN2dfICzKVxsMoWhoXaXLwJDl3XMECrsMTmn8GBLL2UoHFpzkHzcsPlFxY
sBLsw3nfIBDBy/qSlIgQzifhLR0EF1BKNRTAwBrCAGRFUgBLEQPzVk3c/DRk/2NPLI+NjbZ5SmA6
dsqv9xMMshYhKAJNwFqqFK1jBNteEX5Z6K+qls6PjPFjkgJUJt8l7pdwq1euEh8eyxgatWPNM2OP
+9tWA9InpitzpbWxtY8ebvIsd78zquEYzTwEY5zZ+5PjHDNDpSedVTV8ZBm0CyvcvsdUD1K6RVBB
i0fx7bZuJ8yY+kxE9Meb6FNCqoZOF3KxCEfF7TXZH4uL0H+Rv60Iv52+6Qifsh4Qi8ibGXqRj+g/
sHZ7gQ4uXq5/g9KShTrM6w/MBa+4BDY2Z4BpilnO1cFHoiR6DTgNKEeAePsapKWzXyxte/OAqg5g
FpvDpgemT2eSfViLv+NQT5P5OO5SH+kjDlTrbq0cBd6bNK2r+jTBj9b5aWNgxrgdNmo+1Hyo7ejf
rfcgh6SbAXeIeiW2wBLZY4u2gjAOAUpnwBQWBq+PNKeS8nhs9kTqfTxsmWzje4LzvO1hK9N3tXTl
qNTfoNvi5mnzhSIwMtU/ukFC8dCMVgbFUiTzy763B0rjtWXOgRL/NQGcEyeYf7Ret3sF5cbctOdr
05SLP+v7GO/hv6UBiZDJKHwYZ8UuztLhc7dSN4oEOw4HvZ1w3IRqXSqluN5ZJKFoZHJsBGoe9yll
PVmsmT5VCm5xL6L44kRMGLdXxXvIcFIyhLyIIRMoNWM6MS5eQ2j7rJxRi1xA0e2fZx8tqQoi9SpZ
J8bm5TJFbaEAYk7pegvM3/f0G3jDXrXa39FboSSbz1lcAGVfj9JobHFE/l3M6b3c6WaPq74FRYvM
pr0+nDwILc+oezZazJuc3avxv+89DDgsheCwNOmanvRGlD3l/VJV8Yp4/uMN5Qz0nCFgjTZiasZz
46rIdc7CZE1LdKEJyTWD6qEtIyeZBKVwP+cGS4s6Qq7mpRvyhn9vrz5D/7doHi2YP4MUr7YOW1T/
HvXwGhjv68btETgJN//Nw55P4BEIaV2rdozhyMgb/9ZVxq7fX3TLlPWbr17qLhBbqukXlQI9Pxqi
1oltEJrWvrxUOWvp4KysPRrYr6a0kR186XmrGFWUEmbcLpdZt1/sboOznnUNpapw4EYnT14wbO4x
9kUGEf3+O6qPEfBzYQgHNFwRurocrn9g69XUxlml+Fn59P/4uc+K2eABSnz2tidbpTHqEK9q/B0m
El+N3Af2Grwtg4VA99Z5+1VrEAsQUOJB9FE3uit1zYKCwq//QJiMKfOu+MxxEFGWC+EdE1yh/MLd
aK8fE8QEr7xrBQpoIJIjLkgG+/hpeSb8mBxmV6RjuTwiOW2A9llg29nHg6+vVFyXNVHjiQ9hH9BS
WNUCpwb6gtM8QNhC/0NrW13QIeDLqtbK3QzjbLj2/gKOGYzfjKO25w9RAymgkhV9IVz5ne9doIgH
Pw1Ox/uf8AHaurkU+eVN2jASuGOrTmek/Ll6Cz24BK8T0AJEi9sTrzm/f8loheGpNGfUYudSbjTu
QbEXuHgArbb8kxoLwhgBl7p1nDpHEK85CC8SfmGIAB4TG1h4v1tC1kBjsrpBEVJab0XSJQLtEZhD
NX70iDwZg72laz3ipl+A19pJUyPsJg+nagYmtFy10vYWgRABi+EeWhaM/LQE/lH0mVlkq1eLLfct
ZR61POghjh1Y2ivHgooxS4ZeNtsr045XcgSAJ8WmymjZKLbnRrBZ0cQMzhyuGsnro3kG+m12yS/O
OQW68Yyn/hAGGkX+kWwzBwrtD3y1zPQftYr2GGIhrL3iLqH3RrGZ+uzxAS5s1DuCXBjv8aF8yLXi
8QhFLC9T8zkLMKWWnO/9k9Vbi7tbR/7eJwef3NFhkpacGUIo19uS24mm00NGbrwFFqrOZAckOM0o
mOQ2OQIGkfJCnxoADz8gLAytJcefb0IFuzJU2JnZbdZGzX32xmG7zU4FdQ+IFBVOBHqcJNEG9jOB
Y62XiU26AuWlzloxcx4vQ/nN9M4T8vNlGfFLXIrCnwAvI7PGCxjo8sl15XyyCtUGVIaRrygPkFw0
u7k0oBVGFwNMlj9vv35b22qlNTOdGi6hF3tZO9rUwJpoAaI4JlYn6cpbpwag+8UTCmJ0/CPCOJMM
uGNzBFXoU7B7Q4cb/1/y/ZPo+ok3NcKv0GioTZM2KW/uWwiuef74otKlGPFlOaIWGJvEKqCp3w2H
2QlIEbXwN1a9GQ2A3HvHXH1zxBqPMnqNLC2DYU5gvywZ+hZ8xrUcYsXtFWLXmmNtwGydL6h6vACG
GC2zSTPgEr0Warjx7ZhzbDOFHeqvNq3WN3H2rYxDXHogBcUV1/xmWeqfdBLH95CBcWjkzYiEfhOm
/iM4+Aj9U2OhqK0VsS8dzIvXwAkbi+NNrCVAzM2VgdS8ZQJBaYlS3K9fzBH1WjQLr4NGfR2dohIC
eijL67tDAnVzTVXBENgpReRGiYIdtJtBOrJ1s+NrCwFiayQ9g2drn6Ok4wwjEv2jfwUf9s7PRrht
2x5XMxLMFOoGlV4sFxbp2UyW0hec6LVTkn4Nv52HsZUHFDPnhKdeWzCJGzqu3Aa+IrRVRS1X32H0
98pSVhdsglq1zZ0ckDT2IDyFHgIcK1VeGPfZUENw27xQOgUQHmCSMHGnEAuk2qNiailmN89b4HEy
kZi3xEu1U9IAWeT/LQgof2WuhgIynTQgmCkn3QI6ncuw2AX/Z32WLn/gD2mtEgSceVYy0uqrgN3U
LdsgkhqXcCbwFSnNqUJPj9y/gYVoESBG5M76EmptQrPW7iLej7kZWK1JxYZDjW7aFQnpT335BWQP
4t9Dtbld8aniCjYJ3zQ5oFaBowXlUBEzC7mB3llgNa9Wph82RQ/atMFt5EKdY8+jZ6cAS3EH2ITD
upyNvWeZtR3M/YsVNna4pK4zqi9g6ModkLEpXR/03/3Pwd8urVHwQhvbXMwrnxR1KX31iI4Q2Zs+
lFgXtvzowi3kXZwoj2WS39WwhhF3ZPcmNjXJ6t7JfynK9whSzd5+NduVqlV8sQuDlg1ZBTjtiX4b
NfEUqo/X/AepZfBMuoAszc2qPvYo8Kvnib4H0+L9duTZKKm8mb9qnYQdNgycxepfMeWi1ZWzDMx7
YTbphv+lZU3fEasPCGwAK+O4QQMLgvIyJhx61acH/NOOF+nJiTYHNWayaxl61vB8g0p37Jv3Wcpd
eAGCQG8uBVTNORCTTIVnVw7rsjlwLU2iC6vgl/S2E/FikBRweklTSsxAakXiLcVINNKov38nOLp/
iP0W9CJHycm8a9xSrt5kjvMXOL9ZFllIJB+AVvmc6ywqC55dxnvKGqn9Lg4jjLq/O1B+uK49qOy6
7+SgzxfdOMGl6zVZvDSc7z0FjMMOjEPESgPCCn6st4ifqv6zKsjKMj+8l7hUhhXSERPONFmJGfLo
I7mOGJFK/qbZqOdmiusOanq8OFOmmXSg226WQu5kJpmcz7wJyhASeHjp6Sk/+gb+PdmdMQ/Arlem
xwhOQaUMckVK4M/fldXJqOIJDLBYXBqkgmEd9sI5r8T0zMH/sF07djuZLr2HXp+u0a4ytHr2RKls
S6mhsSUa7/xOOoSVU4NYZFbD6T6KeGQUZa7Y0AxD3Zc7i7dx+xUBF52mLvh32BGtm2rOXctoqpay
jccI/YLjV4hLG6wNXnvICdqNBVJE086PhLkiGy5ui4f7nXkRKmnVnLhwFqpkiMbpjBsGww2+xDwk
Q5pl9VDaVDENLoNSGwsK2Ua2YhykqvZXDIovn0i34oVFNkMMSgRxExaxvi0rDI/psapm0JQRIVUF
+WttZdLqN6C5NKOwlqV/+T2U3RBxjt4wUUtUSnH1wRTpuHxhEbqulgeOndoOPSd8a7zsg/30XJbN
bvms+wpK7WjN5MYpMMhA1nwDMtTcRVinWmbu6ljRFA064xwcjAqs0o18RAVUA7YiJ4p73nrmDNy4
/5f9VEFng9p4wmNgv48glGbJDQLbSDSI32YKfY2Q7AbsuxHWOtGx/yWJPkeEeJvTWrUWq1XqLy5/
nLvRPpJ8ZZIZqoipbvDhfhA6twem+EBeifGB8R9VbWef5W5r+HJ1H2Vk/ofbuytY7xVTUlyEM8Ph
0lwD1wgBaF8b2nAhf4QPcDDM8903l8sFbUwBJ5VzS4Xx+WUqB0OTrMr42r5n25B2ijdQuJAZNl5S
Yw/kcC6Y06H93gjqI1gYL/tP1jBXOdvQk7xs4nvSRnI26cAhjbYftBnzt3xaIyN3iDdYS5CUlhQ7
VOPez1YWQMSLj2PdcYMNdhJw2Yq7EOoH+pdQc0DrxQSe11hMsZJCVqwBoNOiCvZTeNGzuzrVNptI
t/shVW/Br8pz23QGvzNRtL3/A8YE5XY8ebbz+7M/59a3Hj+3zmSp2GQUI46Ho66p9eFc6oFS3TZP
fwdOt6nvtOafqT3vmljloFBozIXqDLtmfV3qhxqvC6xmd2WCQIWqDgF2OPoi0/YSQeThIbe6gFjC
R0Y38LEjy7LKWjYPR9rUqFi2CKHf8sDZ93P/yjn4dbyE1FGXSNMmUMZLjCQaa+mF3EKkZaENde/I
7nvkOzVQ2FLTE396mctNvnMTTKecMYplZN0f0YODwPsn1ae+qLtpQim9XsTB2hsTe99Aem5BXhsS
9oqweirlaLFWZ52zCLiW+InUYnVs5O5U3W+7Iu9ZMBNmljqK7KqOdToXhZa2BoQN0wCLzzAz0ejT
tLwAnYKKGtLfi3HD170hrz1TAwn5p9tl6iE9iibfSPG9xTtRvr8W7EcL4uKfgmqEb6aYtbyWbGsZ
7KH94QZhF+cQNZzSN42F5UFhxBL4OjUWdrt3i2XK2ejrX4MwbO0HEY2ZVwn7OgmpItVWgjZlwk4b
tUy6u3caIhJfgfYuzkkytWp7Aw9XNpZvDqk1nl9YS2qU+T7bA1bryupz0PheOpXvy1vgctXluuDV
6WdfnUOniciPk543lfEofznC3a2i+pz2pKAor+263NYQZU2aYBqOr/j0Rc+Z+DChD7kntQOm++Ij
/VNERzxG4f+5PokPkU9jXY4MR0NtSCkX6/zzMZHBQy/wjyCPS1nHwqS0YpqIh9o9xacwsN75Lqtk
89ZnnJMY8GeV75Bc5LUD+HAmtC9d+oTWoIkrq9rdJjXlpc4U2RTdyZKT8S5md6My2f3hDIm3z2w3
rQzDPu0MXybnxk7rrxZfuENNvTijSkr0S1l8L4Sla74RjtQLFQ00gCIkn7foj2nrFbQMX44ERSF+
eVhX2V0zd6XXFIzSHu4lduHMonM6jAnyN5eWaVGKGaVpzmQaWp8o6701qT06ttCAp2pcANZ57TcH
6+pNSD77W7D2DmBcnFdOKc0gE4/q1+GRRk3rGcX0IIopxmpgBypeSuo1BPWP2MSqW8CkEopli7TX
4IcqLZjj2x/d4pP8vAsRkAK8nae5fMM4oN97hPG5hV7iZIQ8v8ud5Z03rw/JT7yHkp39f5xvPl2P
VqexPtyjdU8FF/2+/ibVYuWoBgcqspq/BUfyTqKXBcu7kWA7c8/cA5D/U3WbnlEm5FmLfdAEojXl
b8KibSHzEg5w6LrAqoGugdd74fsHEbFtZniqdWkdNEQHGeAQVS9Lj5j9VElaP8pKQ9zhfzv8uRLv
85saylLZUzX5ref+RisYLChSTyA+eiTOFJzwAb2+6hrZufZEQonUTn8thHgktWUNdLcwVuL3IPX/
KlbXXZlTQapUGJke5s9fyl1sOAyprdW7jRmCViOXX6qGkoqoYNoNwiux+xyu9mqak0E7ITIm48ty
pl2NuAhLxdx2fTDLTjyrGpKdLR5RgqfsezfiwXOcVauCA7s1CUzuFnCMg22kNtopGMAIoeGVwMOs
n37BReQPcKoij2u+usZjUlNoyRo92D9q7aNB2q9mj8iH2qozq8ivcDHf9rw8ZZL3vbse/FrycIcm
imgKFDtEtFbopKlWI/vrQtMsjb/mzYTooyXIt23A8+f/DiLa/CXHaSFycZEd8eQ2JY1ITAB3pJPm
liChDbW/4OnfayWIUFd7m3ZZ/IKLaRQ+cGnf/3514ylNQqiipR/g5vVy20LecNcgkuxlu7QkbaKK
BmGckPw2EnbfZF2yJgdds6eyjH9NFjDmOR9mTfA2X5N67eFOgMNiB9NMBzPEtFz93n7AyK0Mlx2A
m6PR5NwYJexvh3+BiMkTt1eiqeqU7+IHQpvoR1L9cL6mZw83pzleZ7VfTENdARwDYiDzj/tbbmmf
15wznNcuIgr3/dWGfi8aZEnyq56TLC4Oxkp3Q0Cr4ADBi/y85xw12ZumKenSzjI1fL5yzfdUw4tP
PL/DftFLz5baCobM8Uh1SPm20q4Wtxy7kTHKe5oLxfyL0XANqMoSwVkUpBRraCre5kBMJagFXYnO
SgXRwrGYO5j5FUgL0h+fVkonhmetI4B7f0BomDaExB8dNtTcPGQJLZUYwBaQi+8yCrnDT31hzdUe
5TIvau1xyf1eAHLGcWhNoVKZvO4lgxA4u0KXKWXApbV2elkjo2NDIamxD3teaccBslhXBNu1qsKH
ocK+EgBVfAVRre7a+2fUZr1vr0pEsYzQI/iVOJVISCvVZ7TinNeu/1LrRYbA67SPaSq+DqBw9lTJ
iGojCV3lcEAsIemTwDzYWny1LcB55T2nQaBrk3+jAL96nmqOZWAtX40BSsrcQXDLiA5cmqQ5pxIM
EbnIVsD31mG3b0ai4XV43YATnbuu17z4m2ajODn5gGf8KlnrsNIehP5JoBhFFxj9LdEgul3uwh7F
t9ILRx3XGeISwI6nCNjbiIqW1jy/0LAm3G0xMCdWuN7toFA3vDKY9YfPdV+w0glsHzqCYdf79imo
0dl2nwKDZXbDTifl/Gj5vuZNm0V7vdlO7b9BL4PaQ1nQ8igXfjmdLInWRXcA8lD3EInAwcYum8OH
+5Z0gNM/XbWKcii8K0e6B7xEVhr6h6O/SePnoig1cS72crwCEk93h9Z66o6rSPpV+tE/EViAI3xk
Wg7Gplzww4msplFEz2v77f4Ble+s01msqpmVpr2Y48i4Mo4uR9HKWqv0Riw5C49dxlM2LlUgkIS9
1IUFmyHVlpXh+zIliWBRRUlz3F2YjvXViueGJ4/md8xiNz5W2alA2wTsIDt6GWihELj4dwg5A9Sq
sLOT/eC9APVvbWnujKPz9l3ZTBS7wtmMMtKYDZ2oYGCZ3aV/zozcyDIRkTteElcw2AqM0XFAaLCu
VVw1IJVn7VaZqx+A1QiY4Nmd/Ia+aa3n3cCcFrFhk9x4cbcbspp+//jDzkILT0SheNznFknvEJkN
igAh3C6sFCm405SKcWTT2oIzL1y7UWNUBvfWykVUr1Uo91G+0p4btrYe9oMlOtakdUebr1dCl7QK
WUPyyG3YwR1P3jkClGZ3a+kPLhHmnSqOfrPbAGoxW+Ob87EN7XlJrBWArdPacb/B0ewlYZbWfvBh
+gqxE5jK7JWT+rXKU7n4gcXRSHEgf1IxLVfcPSHBUCyWSIrn12Sml/c21tMaetGqJkCLWryEtBxh
VvbClhduOr1HpgDBHm/qojyWdXmN/diyIfKsMJhoTWI+CHsKGhwEYVWNZwQYEbLl/0ntd8LCkb7M
7n5IY0dfCHdQuKf1gyHCoOsfa78PkRYftUYy2R8zU2R5ur4E8Tc/gca0puQ0twl6yo/z06aok3Bm
S9tCAPuYaXJQJh5hF1RPS5kn6Rzdtk2HXgab1J8sq0TyBeFRsxuFDjrNU+WKFhDk6WHwWQAVut5O
QqIqdR9hP9OCTN1xhmaLYUnAViFZqSUQiKYI+buafxPBOfCpc7bJoTCAE/XolZPsxLnE86K8MuDy
w7+LpgxFBZrbbTOpTu6SKmLWZdWpsBN63vyexMFUg3JozdvPrVdptL4mGsynJDm4mddN0HjSv5Xg
6QT+ubia70LVgJTsmCmKEL3DFYoqyuqI2QJROEnyhl1WkhC+Ag1r18d729wAR8Z9nwyohtMpIk1K
qMICPm3xBu8G05OB3TBQEM5ok264+hVRDZZW48VZAQ8Xf//VlsgfBwsRhS0948kN5vD7wORUTdl2
9+5PE0u4IFl1ls5PSlhWLWr8boSWL0DERQGmnVjA4021d6hGG9PkRQ0rvb01aqVHNyQCiTfdEE7i
KRQLpHyHyMsIhOhC3SVn8zid3y3p8opiSpVfsrDpc20oO7X4hSn5+uKP/28SIC3z7R2yxt77Tgkf
+XuQfw4PnA1cPLnRZFs1cV1jLdQIb11BlsLLpofw/Ias2ffiLZhIkmXZXlNrB8WoWkEN0SNkDuAE
8WU+eFkcltuPnC9Kebc4suFOakqF0RuF4mScZbCiMgqGXKZGcRRDrMZKLeAEj0iu89YuwgIitkxu
kdgU0nS6h1tScp02HLL+k2J08rR14TUC3muAcQleETL6GAvkLKzGuTrK+DqaaehmK1j9Hgc6JGau
rYKl/l73INKgDKqE/Brky2dNFkRBVjVEV/cCiUndMYf5wWO1odSpcj8JUQZcYpnRLz8rYmU+C8Gn
SKbbnbGXHqkFbs2WH2nQes7zavyULDdX3W4LABOPXoZoZCVo3ZEuBanAu6YoxgOkDArwruF6xran
2q7+5iU2dUb5OPQsYbmSFiUwSxXFUY+U8ywjV6mPQ/DNIQSZGWnlB8UFWQOmsJ7IsT2J2U09aa2o
+QOBat/K7ClPgnIZgykT+yIooen4YtuIJx+zWIvHqEoB/hrAJ3V8B5csNIdBSijRyGFg68OhdaWl
rNxaI/YLGjG4sn/q/9Hn2kMAE9WSUq9CVN06UJdcVBoi6HQlwWvOOrmxTnqCaLIUdsp8NbfcXPHx
7YAYyZEZjTvrbHrCJNxXqcDYBJkGa7SHBnESrruHXAlSUNyCS3vnGfSsC1FWoWDV8ymzf0U9Pf8c
zNDkwP4RqLmJv4xOELjwiQtvQrDgj0btzlFUlgJh/mGII2865gwrIVDlPMDY067NJtbT2j1KEJeD
QS5B0ZZdNVS9RGInPlcuXmzFvo3++wEZ2tPI12mZVd10gzIqG2S3ZmZutxxcvczXK7WjIRsFaYV7
rUI70zUJkn1eV97uqd3SckTkC6utGgeHkzSGr0w9nlhJJdrO6xvYQDEg/jke52MAKt2blJI8HRjO
Kksn3zPUOcxvyACJpR/IkC/EffX/3t3PHkkR4axfTpYB3LgAvWmeT3aJH8RKwYJoLRfmDtoQfH0i
Pd3k37Y3thoqeHNdmcU5rRnXO0nFqp933Y5XM4m26VpPvXZAeZ9LjYPe/dQBel4IHI5+UqqLZwZT
JY8NFm3vdrOKy+I6YPLx6S2r4HaqBgFIZAqzYEmh1BegAU8HiKuKV+Dpvk0NkOUiXtwT+ohLguf7
mpAV27jh1i8Lq0roNkMQ2F5lDzfRw+/KIFonH0U5HJiKELj7H9AcBLTE9W/3ZLIlTcoRf20Qx2bX
y0kmv2F/LnZ07A6pwPjHIJ+lbmaoOQxrZB85ch7zdpU7M9YKjndCKvxx7hal9PphZ/FAEVAsazv8
8i8143smNm6IlSbBohj1EEu8RlRNGk2jNer2zPQIKOHVBnJucNcy0i9gUaUTEkpaTih7poK8/vsp
bAV/O3sqUwalL+oXWih3qqlQhdM4pMP1RPaBleO2JfKKDOvZYG4OrPqLF0IeVtHuElvsIw4LXwn4
4WyO9VGi9WQE8348xmo+nA0wi8JhWIEKRAtALFmxdP5mLCE6zMe4b32X5Q83z8lgc7qImuO/9zHH
MWP28GzOxR+vmoszQ5H2VEK7jWkDD9DKaq5pdNComoGHoq5Ba+8Y0ZVyplGY9EXbmf/fDg6A7Jv0
+NxYA830Xbl+PKGPpv1OZAez1cS1Bl+NehP1AcZEUGFfyxbtoi1WYlOrokyo7fqnuSRH8culUNLH
7gCPHwYqODegrA/zn8YnTjLTheDtfKtsGI37EJ5MT1ndRBVT4KX/17xnZXlzZaIWXjz3JBOICGQ5
ouJu2kb31AR7iwhP1KuiShFKvpCo3AYQIGn3BawvVgh1PGYulJhWmhnM1AtliFiWkx3h57fOMvyw
L0u/gJ+NEuFBhGZ1OUzoCTTQEiaC+cXS9llX5iFLpyWUjhvuGNCTwZGMpwnbhkfa1ZjPNmtHETGB
i0P/xRyZWGFdNwvf27HMKSZVxoErElJDgSK5MxwqUvOZOiM/uk8pkWRaa8g5186+C+q/ss4kekVx
zxTIBAY6+bUmLU2g/vSyX88ZmvCz5QfyoJ5hgnpcHkMM/5hB/pqpQBWnylEbeZ8S0wgO6LX9UXYP
OPmb7Bly+hYn5CKr6MCgn386LUbl/WYdqmgLrdQNLBJbcFR619wkrJU/dVInS6aKr8HvzQkDEgdi
CsleKr/qW/KfflYn75UGCweWopLJ7KdR8PrPyYMPMzotGD1gtQBEal/TqmWkvvEFszPprF4xwUpP
mNYqDjFBozqG1ond3fRYZ0BbX0eCi6SbpNywZiGCB8XMHNds3PfHyBhFUsh9yP6Y3C26wfHsLFWY
s6UAIdZZlXdzj9bKax9RTTsLCY0lfHzFWhiAbhAKcnhPqf5jM2WJZX0MyiEoLBBcOeh/a66SAbVo
n7NzFZ5GMrdIGJDOkqxSSgZdeuIIzi4BLm9JODcWfJHGwDDUdxlISkBpXp2uG1SWEZMpyF0/+0Hn
TX8c8xlMbs5Ga4CTPmOzaPBQY/LtaBK1Sqv7FAl3II+hYJa626hMcaEoQnrXTH6KOvu48aT9G5at
KCviW1xW4j4JxZkl8idTtMZHnOuECTTSxmkOQT4azcafQx61X4gc0OBFLSzoXAqdWQl70YhJb+J4
MNLeU4E5BxrwemDk5CFqzD635up+sdxILC1Ym7gMjgRbo1/G52WfGj2rV9PXQ5dFAxdpyMQi61Ww
k0HwJezp0rpt3YQ34iR/zW15Y3wg3nYN66yQylrefedL2bcWxGMZzN05un5sbvtKhBjal9MXN971
ZQg5SHedhzLAO8lzP6C207JZa64bA+LzwevlHt9ZG6Oa0DMV8+zAUroq3ulRfBlpzvPPLoRLJjVB
GOa9PCWzMC9oJXIfL4iOk1g2fQtczmhA9QEjfyxCqMw+8FVgsqZp1IEoAc+8uhafgGHJYp1KeIVG
IaayuR09nebsl4IdpgbZy5+CKi1EZ5Pp/8JAX9FeuNPAwcRzPeSoOoxts7L0zko9TsIZzJaKSdny
M6gcb8MSmGSITMRlU2+8olGg5kuN7ODthOW3qwtTj9/6rL7wY6dukzhxWeEUTjZT/Tucyw3zdhKo
Gd/JVe8paX2Lxgu51aBxZAVTej7NRdpKTk0NOFO+wQBVbVr6eq5ykQl2MocipcQDxkbuC3JsscX8
P+OxKH8sl7YDwrXfepmGYf3oWQEa2YlAkbqIWYuSq4LtMBySMtCEFOWKtFTNXR12SBXS6e2VqEm/
1PYmJ7F4vw0ZcclcZdQ16Ev5pJbKyqJ9dGg38PteWUnLv1YPqL4gELv5MABV9jN6tfDUf2pVtUBY
Ysb4RN+Vb0m6Nbgac20Or19+2YiDg3KVnDqjKuqQBmoJl38p5Icll3jZpJQSXMEDn3dFln8jKJr3
3mS+7mOUrPmzf1fu0LpGHmP4EjQqDU2mTbR3bWG2F1Zyqu4o7UXw/WHPhcmyzCw48SAF5b1NQ2EG
jUbcglwqvnAhQyPNPUIiMKWxf5GduxYM4ugGG24z0pR4//TeORpoee1hjtkIYnGsmRsOcLeOiD5K
EWxc+mFJyEPT3gWxG8pm2PsHALGzGiYevxHtII3h7ZEKDEq5QT1ZUkcOzMlZFL58ZYgQeAzM5YIt
TEcyjc5NV1JU9U0QCIayn42x20BmMKAnqdjugOJkGpHUh9WYhT2U92ypuWt+1rsuuSIQCyeczWlQ
SkVXfn7XmaiWoyPdwpHzU8OJ1Ivx+IZ8/X4w6LF+d09mC6OOl2Kg9+ldjQrRxXAmcap+e/ulVz8A
aEz/B1uAD5atnoh7+rW+ozwxvbV1YErRGe/EPETT8DZu7Z9vnQAhdKbMFWVHjka2bHhat4umcvfx
ig59rPKi39/ZPDe9P7hNRK7wC2qw4p/Qp0jeJd19dSOa/bLVQta5VVxcPB6KAxFkWhfB3otINl3W
uT3ElM75ZobISwFYv3PvUS6nadrIIasLmK6kBWpG2zLX2aJi6lf1i3QHfYuFTbArurkmGP8CSRIH
/xzt1aRQ3rqVCzkL3qv437d9tmUD+YXOqcsGK9ynihwddxwC8Lp1hxBnv+pex1z4oM+r9i+99Y7q
M1JkJFdICWXH89iQoqACWVn+ANWd1p20i+ELyj9lpl4FCHfYDIk/ZGpSilNVQjluWAvsRzqKDGns
hxAtFOEuayGT+fkNoTggMx4slcfN0P4OQ10CcXGmyAFKGTdd8NrQCREeIFxgZkY00G2m0DAgsLsA
0iDXxa2UALphvSePoYnXcSsLOzUI8TCCDC8hIg8vMoJXX1IO8aJQ6zYc5R0DLrzzg5lMZQCEPYyL
CKkgdG5S0zDawl52mqh/JRUDjBwhqP8J6myCQAde9xDLKpQ9GHyn9pg1OzYoID0zEI8tyyRbSJem
1TJcL77vktGe1eMIhVMDSACPMWxmBR4Y/wmd2/xy/p46RqhvEw4KEkPahwY8CIEwCvG7QH6oCGMU
XMB/v6jyPzNSWnlMFxxuwOLpCS21S9jOUo86HvOG9bbkSPAS+a7C/CXg49pAP/3uU0p5v2yz3P7z
/kdDOzCNVixkMvP/DW4HwqJU91wbWi9DUPN99Yhy8zryrmWbndAve6YXWcSdX73P+Z3u0LRJd9pH
IQIDgieYBSMvhs2srjc4DQzuJZ46fZt5s5US4hG6NxdEk2gVQPhkwN8F7IaxPK5fvPdEA8kTDQ+I
gXL0IayurbcWU+YuTue557mCqIwtRypBT3h8WxBKuErvg8sR93SX6zrykteW9oESNpIyGy3pYxn3
1DnKhkh25rzk8HLfpTJmcqIsSTCVne9EcZj6RsSQLpiuACZbkngj/5pNzImwkUIrVixJDG3xJ8HS
0kbWkK42WYCFoU0yhNSRXsyX7mdkKqgpMQIsag5QqQJA2JOEQPn+LRPXYCoA3z7JxFHS9tgXpTVL
e9NGCRm2C5oEnKPrUKxTvfKGCHOMAhzCuus5qlm1YSMLxc/IIjMpGPiHOUqU8q/7ELXn1GaE207t
Q2YQlC1H12u1UYWYZ9oxCdTiyvID7wK0oe1vskp9aTC9HY5IRkApJ9lYikupZjVA1JtzYfZLbDmM
Y4RdOU6/G+Znvn/1B1+t9BXdH8FuP7fosJk3vIMdunHSltXqiTseZqEybLau/b96Mxac4Nkq+LbH
H9Cz18uwJfhKTDZjuZoRxZN+4+UYE1EDxIOxjiShex6GftP6/VRyz/cm5sYR215blvNA9I15MW+o
dNkBd9739yvJsEHfh0UutnlNl8Wh5i4nR7nfj5ULTln01nhpVvOAlqrpPVNpDxsaWsJSbWa/x9Xh
qe8j2HAgOmBBAyp5LAOFVHFU4sjHSes4lxrfVMw/2iwo26Rlr5br0gq3QSD81Z8WRMp784OgpDmg
2OJIGxNdPH+PYvRBQJmDejoRB6jO7QiOvxdZk+3bfBnHCWEjWvJ+7RIA2AYxVZW9fx6vKnMt/wMP
3jc9AKaN58fVjECUQh3Cjd2md8wTewEUIVMF6/GRwfD6g+L6gQNUJ2ZHgYEhmePAcBGvo4XAetgH
cH1B5Y0QMy15jOls+JQ+c/POFllMj69amkOWaA/mmmxWkuuJ7ANJL7K3ROa/ZUgRw+U1mCYr3x4y
Nl7CiBoRe6q+9SWMSAkSJnDKl3o+Yzdl8gEWjL8tA7vZrQX2QW13XzyMU1xZtUMnG1m7WUrYnuhl
jYWSax8gvbxjEw6I0f+900dodwA+TGmAqsifHxNL7oEsxiuc38V2BUM1g/z3qq2FmrKbE3nXuofq
ygaYJqbhJrH2E3iAZmkLAmSWMAn/DoBdIK7t6KAkBiW4Hi5lITTt/VjS+DdaD4AP7qnOduKLVZEZ
/x4I3EzJ9dRaqU3+5cDT9RwQDiJfSfOLn7aAueBoO2nmFmTVUTkjZwU1gRG3dQgYwP7C4YManI0+
CZi78aApp/ZMaZ/3mprdVlFb+yCRq6HaVzhXjRlnGppy/KiTe+2glWfiaY3TvgyHgVRh/N9jgt3/
0UZlenwUHDLDwRv9mGlcVWDTR0J0HpACpWowwZEfap84IC0NwW3phICal8DVa9c5TPd1hycNXUFI
8TpwC3KYVY71zeV98NQSLqdRbhCfHIDdNcF+hLC9tNWdnOoZ3Ipt3BnPIuSUGniKQT7VRDeDxT+Y
fwRl0n4dS6RSk2hFCr51HTcDhqnv/YgUmH/ji7vQ5pgwnGyir0FZVRkYutQ4Vzew9lz/PtdTwEOk
LCloswt5oQJCWnz8LCcB2qyeiHt1eK0+owg7yUjP5OMRMcH7NPRqjJjHrVuOpWRnDHYWBC231pXf
2mujXibr/4e2FkaXfYUTPJlKx9XtE7BleLOKrpSefjZuhf7/mKqiG5gjhi4vchTEhJG6JFVRGGMz
swWKWQdNhVnU5WjZCVbD0yA75AJedryKbce1JhSkWGa33ICuY9Qaonn3oQ29MEtZRsVqxZiBtlYu
NV5RDAI20ZjQImu8E8gHpFBTun+hPPm2SbV0duJHGb1O8MmmYOZpkPhrzLO/3zsL2CMOB/9+R+U0
BavvyZdL03jdpH/W5TA7v1IFjEUkRjEuYFGFGldhf8wOU7qbEs+p3+JMYqmCW77Ml6bCeb0S79Xj
HTc2Sejv8A0FbN3vBZe55WL963LzAdeyNzFpMklORXraV2Jf/p/KPnxkycbVbMdxPBsY5TuOt3cv
smoVfYKVDh5Mrif1nDPPPTN19Rj6DUImaM08AEb3m3G4ZrrHelrGPZx5rWFIsYL2Z633ZILQ0dx3
RyJJC/ZRmdSzhNER1HM2A/vGVdUe4TGVc7aBWXz7/So1I8bEguMwObhHl9aP4y4funqqQYpQqgap
FAv3JNTlm3ByY3nreF0y42FR4RpQUBEm7+qdJgL+lKoKw9KOGZOExOilpveYguegvOZdVVWif0SQ
rdHz5/W7SdF2PQMDJDIrxK8jJsSw6Um2p7hnUUaFlG7LenLYp/6LCrn0l1ILNFg7GpoPhA+UlrTQ
QlVknR1AZJu0gepmGD6R7TYzmml1jwn0rZvXXD0Kny2TLBRPzCfsF6OepizhjuPCFt4GMRuc1NqU
gYnHAcxIi+uP2sP8hR73AT3jCvRbs86dwtc4hKandAUYsMRG5BMrmmTkGocZblfUpSKzh5eVomAY
SxeoxOVLjJ+jrYJuPAbnqmzmONsoXNUbSTzPLBtRNAHxRu6/19LZkjYwq5HwBKxXvd3V4Ef7EEyb
9zY4UQW/CeKh1GsoGdl1+nTYYztgkZlMydyC2HL0CLWcUqKwh6DTCX43k8oVKcHllnGaDsPWN2Zo
QBLDEul+OISZHFeXkWtcr5M7vGa3p/OTKOBj/QOk7YUtxvz8Lg1mHQghzzkWl52hkg0lzJEj8NO3
GpwtKBWsjljvlwEpzbLkwf/JztK8RNKJwZwB/HcPRyvuwAg9mL1za/hYS7mAvrDjAe+Teb1V5kAC
VUW41HEdrKOuXfwEneiEq5vkMD+AtLgKIgcWmc5MmJGaGih4uXqiGAT3oxUfZbV5bBf7zJdlldmC
mHbN2AkNPiSfNFXJqzSNSopPznvu+SKr623zXCiohnE3z3MuBMtFmNmpuFW1yz5VPks/hrwQHjnV
NchoCGCreBD2l2nqEJOGQU7hKjhX8g2iyMPDyUXRGHbYuZ5ks4aUG0Rs2flXMbsz5E7li2w+L8oa
DoHhCXibMrRCrj2HInLtubGSGAQbNzLDr6iR5uCxxhPpJCpCbquCKc0/TRXlUzbjJyIDq1tepccW
129rNS7bDRw5UN6tThN2zkUoJJqTSkSw/6JB0HWYiR+gEf0GizTi6ta2SCntqP9wHlTeMyYOrveQ
CESoOTx29Tk33jXa5N9BPwdRydTgWV8PVNXIjNtSK2mM+fL0exv3s5XLPHtkrMegX9MO9k6Gt9Vm
vthU8/kjQkTLsibO3qT2SoR/7xvhPeb3R1vypcLTy5jaPkgcJKv6N55AQudkel+CVPWakZXX8Vim
OCbnqgNeWpt8MqOUlMjeipX5A+gnkSQndLqMz+A/n8TLwgbdZ6CKZUT51uPAmLZSYnq5MntSjled
W56a+0qJQ86N/2zI961lmNMqaA9avX9XMpS78ceygrBFFe3C9QuCAI6PgtZQ+eyEO8oNnXcaZ2yq
8ZmiNGwWe/d8LBmLYWjIzv+5Z/LYXgW3R4TMkjBySYwL1mYyeyljXe08HaK2bkgcQFaY52GvSn5A
vPILuzHnbdEDUXX/LUyyFNOiQsPBsFm+rBBruwzUhpDtCoeoH0WBUddIMP+tbTvgaesQMWmOPG8m
LTCaWg4PTt9SCkmTfO0BD4YC+LF3M7oe2CnvmIrs1Om8WrxLSPWwoILI/tTFLyCb1GdzKMjguAXt
FvnZajVWR+a393mjBiuxrjlhrKoFSNTgLAE+1NhZQGbQ1x8MgPpuFaq7ghQygB/UEuEO1ccTnajp
ZhQEi2yvnwNfnLOSPg6mH6lCfXfzETzROlG4WZY1OwaE7kz8bvNqx7VJGyzNtLO/8sJ0oxZ/IQu4
Hv3lEomoRN1jPq7YjXSlEW4zpW4HsEgYrnvylyO3xMIGsLCSN/ixSPdcvh78wZ9vQwh1MBBsYHFU
VgSVaU3IeYWNw5PrxnzmwUjHkwfEBEuvde9RAkztKEPOV7bXqlZ2+IwAg9fgPovPQniMubWjidTa
9KaG3MI3B48dHb/ce9KMLId0gEa3jn98xIV1fuQh1BYru/bWYaFl9eVQCay/mzxMT+zSjAdK9UcI
CSg2MNy0BHUS/aZ8vHbg87mPAVJIqN6Wre+jluOWoxeve8qv/Go3N4abddbOWCXlY3xD7jwq5IlE
FkSpcvwa5bGQ7a3f2Q9HNgi4AMPRQFPuBi8fif15hf/Of8HbfZP2Gf7y1TRi1CEnNpTrcba6GbaM
BSQAE5ESXDVVrkHpwe3COiZq7mb2F52sYL7vXW9kfsCEMR9Zgft6gmgKBu5qzNv5XmpWzIM2f0UV
C0BT6yHgITz37aNtzGxtOQpIzK5hs2/+/hBi2WNl9C19sFl2HMGKsYlwwpdBxAE9A8AR6mtQA0Py
2q461DanfDF9mrboWbPPErYWMi7c7tA8ff8vFtq+Vt3SROh2JkiNx4EWOF8mbtONVt29A9LpCBQX
AnKv5XUgnx14eS61ZKXQq+2AHgF4VgCwlCyRJFsYhMIcpmQl1/V+FrmV00l6ozWx1Rrc07kfp3l1
ie5Wf6XFcXLIAqFkDk1qUJKBx6BgCgFymGFGdw1f4dVAe6AqidhWwCpLvEpGlVVfo6GeTAs9Ohcb
uDj87tOmtjG3/bIZpSibYCyB+pgq+VE/sW5uE3V593LKlg4SXswl29Qr/Z0pxkhrCoQD/KzCLM3O
gZWLaTqKhsFjd8OtBBwkhBJhyPtMC+UjfzIEs5Ub3oracuJLkPXVR/zW+BANkfvT0d+y6C/NoLGc
gZrkuiC4aMiG73jDefjyGE/CKUEKgpJj75VXuZH0zKED8gfokQXT3ziLvS6g1OUIfNIoL+NTmNcl
/V1Zp2MlWJ9KJAkCqYsZiK7ZDTk9dfmxYut55o8Rus6J6hgaEU97TC7NPCMXU2yvMNr7H/UPuzc1
Dg2AStXYbOYxhg0vPYkB3jFW3esvYsUCah3CEkTGp37g/LM6VFR7Acp3dHtok5KwV0hB1XzSdcwI
c7lJNzjAdjv/TfYxpdm7u1JS+yfX+9CJc6WTMOCseJXXqd48JTO4f6ZK4jWBFoCWHzbHyV8+fa7k
Y4yk+/992M7kB0xl2jRkNhdEMOJIWS4IXYZsOWYB0VRChXvSy9fDTKNL6Vn3xbC99j+hooJ4sl6h
9h1G78uNGN9+zPimDsDZ+AkCrH3It2xytrI9G8kHmwbPcYv0J3Ph6erMy1+u+vZm2yLC4iIKAX8c
agaCizrpczZNvWUYGG6p283Kshdb+oH6Gv0KI5nnkNPQJrR7MPQtf0THy0av9V7Hzddy8RWE6Q5c
RrVI38Ohoc1kzi3HwL3eQ8Wxou+xCanK4XLvUXTVOO6nUyjrnpLZbO/FLueql1d9EslsCes70xUl
B2rdrN3SRY9SBmKwmh5rgXbJzb/C1hpOdRuk/U8rA/BpKB3C5eJFG1k3M9m19q9wncwihnV1U8yo
P4WMPLfQ0mCfV8mGZnAgTYqSdYZ2vyHj3Co9YPN0Dy+LZHQ4kHg3YbM3BuWXlPUIjyiziPjXqb1W
PYm8yIHkXIt6jYvsCg5K+aS9x2xs3V6nKXVClX2fkihBqE05gy0mZP8AcrDBIiFoUCfrEgH/oj9a
xJuGtw563FkkCRpWKw7Syr2sZDgGnQqoZbqRm327UdEi8z3U4GKxDBpev01909mcrPAaBn1UzQOS
XICcpxCE+ltgZITwwfv0UPC3pXU2vnVFM6nZDx+iaiozSFeTKGCDSFSB8ATjL5p94Q0c6eJhtorE
+47+m/Oj1mqJcQBbB7QAw/ff+BxbWoirty5OJVmoF1zUu3m4TE3jy1HA2kDddejHblcRs3lB0VFi
PZ5r8a7lPeMUAjHLNP+tH7cWa2/hlVIXwDzlvRbQWuekLTtR3Xbo4aeDaS2VcdLGWfNb7cN7kv3A
LQp7eKud7NsRVtdp0+nvxB2CdKVDECo9qzzudu+RN0JsTN1YVPx+HU1Hp4URkmehph02kYF1pVpc
KpIRjm99Kqs7RfNklv1EBBV1ViQs7qplntVjQhCa+PgB/9U2cDaVShT5+MYp5t99IvwAHfgPUjTk
6PVyEU4TeIfkcOFG3C6lk6ibak6Q0t58vSZh6DNKIXg876RnxiQtfKiHSP4FEWFw8+sZbKPap4Ba
U7qEgSrcQ+o0Qje3RBkHMzFn0dHw00vm/BLhUwdg5Awq2CMaPAy5dg02EVeVaVO/kIyPpLDkViLP
zSeAcsUyqKR+F4DI6qCkBzCata0SzThS/RFP3+Ic7YT2Cf1LzsX5Yx7cVm2+/I6dC4C+tYgKUXnG
BKQY9HHU1s6dbQVS9bS7ww6f9I4H64PjuN91hBuIS5pPIf/OIWb8BEa4dLjHRc4uqeexaOisdRvR
0JX5AIt9jIshwgmLBM7ww16Sz4yWL19oZzJbptDP40dvCpeOR+wsfQcsCOI7NKYpvpIa55JkMIes
dRTze3FB3idIRhjfjUCnmgATsa1J3901FiRkXq8q2/OhJcf5GrrDzx+RM4WjsGxtIm3icz88mYSV
FiugG3IbrBoQ+NbWQEJd+friUJcOYjLoPPTlp3IReJaiUFkMHFKHKNapwMSnHHk8ysFu4gmkK4PI
tzuY2VV5JTQrWyXZAgAv6fo2s3dnDLDIUYSAFQB6d9YhnwKY0vClHICJ8xfMWdbMc9SOcTOsKD00
WLtwd5LRoEcpqI8n8Bhee1xq73A//9nd9h3S6JvnP5F/OCMssONFgSBPwyadIe3OB4GSKB0BD2bl
wdsv6ugKHPCoRNWOld87vrR5rNKgLnBHwmIa9b6gaVkgUXFskdox1zUTBEAvbKR9foZ8CMQ1240m
tTWILQ2vF/Y4zoPCsjZPJev3y/NYw6KaHMwedfxjbbaMaOx7kEjYNzXDSHF0zKDBdhmKBNIlroev
UhEq4wdk7n95aenAD1X56ooyyn3KcLc+kpzaUZ7zn/IfKFDj2rX5nzJsS6yBKSiZvzOG2kgmNc7B
pNCj6MSEVlVbQC/zVPjMh4BwKk7ppXa4MLVsL9gaRMzaiSybRVUKUU41pK7N6VzNBvM2FNwnaNhq
WMYxdpUcfpKfkrhpm2qnqCUCcvFSlStNQzxoZQ7uN9JduBMh5y84UeZoR+98Ozlu09ESnV7xLWcK
76wl+rszWloF/gnyRNwxm64asjKN1Z+8ZV1Pdlc+VBOQZv8baVfw9xkCEMZl2inx8Y9PGxwgsZpC
MV9yhKAmmkyOmF4LQcWiWrrEIxIBIQOLsHRfuJlDG8zffQrXKztq2AVd2CXuy+AwkwuOtUg851zj
5ZSvM093Qr++8T0pHbLYD+GEcQKlbYD7Uu2Pm9MxBqhU7x1X14llDUDNbOSTtd1Mxg7bRAWpGMlz
ShVEFD3X5V653//whd6qara9dPVLw7TSAlPI9anWEFA37bd2fhMnERi7pY15DP7tq75eqt55VOQG
SCPA9IwWKEcKwoe5EutMp+WoLDsOgfUmHhrvjPbuWvltsqtblJJX1jRmEzGAADq1IDrpJyCkVRsA
48/ayRL71FEllryaRbuL5dAYQxF67I46Zo3lLAVGPrih++5zvbsxOy08uyW+6mh9PeiiJiOxetPE
GDJ9GqK0Uyi/dwErkDh8eBHr0bjeiuY+pSfsbAH5R1o4PqmgkCa5o8TX9bQ4ScuVduqqG1w0+Fl4
TaYyZ3tgBdD0lcoKDqkL7Wsznbi34VBhckBpIGnqZxvhcgsq8ncmDkEoOhWscx5po6BCvM/1w2Wu
yUKMb9ljqhiPgBts8I5tfqbhEd0XRtUhO3TsyIgKOmzVYcydv2lCP6+veFUaYB+lhEv2B7On9q/9
YQFnS7bsvcu6xobavM/am+P1/OdfAt8giRVYmMgz0mspZMuD59aXVVtM9wVWA4Hsx794EsnPYhKm
goD+MtlDMCkFL3HaI43bcu6t728w1fVzvKqaDHBIrT7d8UPaW6mu/9VwFSnmZ49F25TbcVZJoSuQ
PfYzaWRA6+S7JN7JGt2slX1Co8jLJWShvTBmkKCUy929l+CqFP3gvS7KyKsM3JRqdzTgQ1I0kRp+
4W41CTbtfG4dkuBn6bQfkoOhwUir/A9y2th6VIwx7nxVh6d6aXgx3UjOJLWQ8tV9RT7odNJ/zC2O
N5kbKcKjspwVjF0LBhRJlZyWwWBVhi1gZNSeNpQmqOrrqsQJd9vs8QEMi6ho3q7dz1JdS6NpTWNR
h+L0MUy4UTJEldy3H5dC5pq8V9gM3Y2fUpwbF7nYFsKoWNgs5H5bz/7LzLaJE16z/21n3HaTr7Cm
5Hi9MsPsmSZwcI/QYZjBqs8WqpSm88noDVfwtaWF3PPjQ/eI0yL8s+ULMozgwUJfBQeZmaHLTqpV
WOdBNemSKRBvpZzhwNFZu9ieNQI+NrV+C9IcoAsdK7pNkMdIbQgNaAAjHpUjz1XShWoYLJ8vzEH2
38kSuv+CvyeAguGxIn12UtQjcLFcXeQ7AjVrETFxh0LiQ+BMLM7TOYmHAP8tyAY3uR5J/VYzUFki
5mYV3dfkzakRbMUYmCJCEE05PAY8Ti/DgNv5Ll6J108FExMxqQbQ4Y681fmYKGphg6TDffqk6KV5
TNNk2CQyrhn5NdlmaWoLl6VlbJomWcDd96i59sHMYa3IsbvOpIlqM8DE5bJVO7m1v4i0BdQjwpjO
wL9bmU/1jHAKxNTt+OKEmXqHiekyyae1YIa0MY/vQJNMT4DaOfwGbdY5jBxvfQtQoXWPkFXSACrV
+kvRdA4v3/PlEy2Q7HUV4IS1bqijU9R1VgMCQbUr96vmr2iG9QSYQ1lJOL7fJbDMa6ZDoifyrtnI
lJ1hczNdOjSycNxSl/b+9CIC+KTxmnlOmF6B+bKmzIRE2ynPNOSa1ufnlvgsXgG4x2PabV7jkh/L
xcVcjOSfwa2Ru6NjL6ZLs68Xs24+ZZnWOHpzP89haPVLHrqMxMaP+G+bf36RJbV1T7f8o9BtvgbH
0KqBPmIOTjZeLdY0BaME8IOdOb8+ZoVzjo61xFROiJKlcWN/HQoUZdpCkMMAP3AOkvh84u8wdOne
mwtMiJM0r52uug5fhpdGin9iaZTEnuALtM8gH4wyuqhggtAyG/h6KkoeWtpJys4KqEXiMeghfygt
eRRZz39Px14TAzbiWdnpDLM0AXaHWfD4qa8zDyv7BaZQ1yOE4nO7Org0f16XOIJiXJxpAy5rzZ6z
Q592iGFdFH0+S0xDzQvPghOfETEOcgdP/rkFrYDMll6IGtdgAmzyKLdLIi52bKexNbKAMyB+EoLe
Nnglds5jGQMcsS6xsJ1HpMv7z52zKeba/X65yCucWFqEs/t1cdJLNMytjJdmKfChXB/Hv0ogzq0J
8Ghr+0/BkcSFNncA2zAYYdF+cSPxhXYrBAXbED648fZb8F91Z/VyjPD2o+30cZhoXOSzhXczykfm
o5RRSUKKUVM8F8ebn0KB5ibQqTAf4C9AgKiAbIdqfweuvutvqGoMt9j7WziEKgEcU5Fw4yZBD0W3
tDJKZ0RmJCK5DDKRfiLbeYoasqXMfSpxhdHML/lClw973qdfFmYRhRh97TBcs/E3j+6hS1nRin+/
tnEEL4mqLCfebx6LsQ4fJouUfcna+S1lJXiMNixJfraWw16M4XF2tn5X2/KId6CvlHonYqQ1VllE
HN2yYE1QDlyv/uPej9mF8avoYblLtshnvia0f1wKMIHcdPsXnYn+hqHPdJFURK4rmFQeyJ8e5krX
hvtNWrfcfdLPxWftGqZkdY2f5zz3P+HSLu66FxM9txLuHLZRfUE2Pk/QOhpoVKkIeWLwvOyKF45k
tUaCUwx8BMrO+/RHv11SnzcE5W7yO3cCtN68TsnWFcGvdI9wLwuJEYhW1fNhU/2arKvQz33IQGei
NSabepHt0ifZFnE1nj3XrhtWRTssZ2Afkh2u/SMEOaamIK/dz6DxcUxW8X4UAhR5shTLdnvNyuXF
Fz8kjG6+5Tm/c4evmdiVkr7Ih/q6gFNFRzpiyatyCY5ygmKRKJdN88tejD9RmQnI9GWTPTUGca+f
ZpYPrsJWSuoHnMaRR7cvEXthCMQKflZesyrcllcmL6TBb6qizbFy949Yt6SHNJz3Q7g7BlbyGixL
jzpX6NYXu9atkIQpxv+lj9f/qe64R0TnJuKGczeb8tdJNoUpvLgVaAUg3QFTeUj2jY1Vz96Vj0eZ
ah0lLmIrByTBSJGVnvZklBK7mwIdNufqx5ptnBD3MImvp0O1RPfsI/ukZDqwxcwbcv7lP+Co/IBe
4akpe11WhI/Xp05HDe93wSlL0zis6FriI8N3aduaSDlhC9K9J9EE7ITXK6txSIFiVfmVaii1tbgw
FAxUztjPzMuRQO74v0DouztKE0kLmsLgXroiVrxP8i0rRMDo2tQB3ybomk7ihnpSgQ2Ov3KZaex6
LspCDztJRtQBNm+XR5pvI/V2AssoLlvPzOcfohpGW9uL+YBUNLt3Iwh7kt2q6cOt/4C9/9rjOpNR
2c/9kN3tIBdgA2ARLNABd5b63zL2n93i5FiNit8g8pqplFSkD/uSVV+/TJg4riS/VajDN75alzpL
Z47XRl45d5Kzbag5cLOaFopnYjBVnLjPc2HATwHEUSvVFSuCnYvnE9LguI7mu5s2W/evSSXZtH4m
I28ehEfwfqf4MZfQwcwBMtK71+GcwQMk6fjc9bYkGgqSndrTazkzmIg3nMPMsbPtfreQcIJXUxcD
Crf7OXJhcvpCOKfoNXgZXeH7Ye7Ks7DJqyWqFm4xbigXdu2FyF1HkywpKDCxCCVw0+eICzg+xmcd
NbpQgf8YhPWBBnwXhqRij7B/E0Hj2kAVDk69rNBJ34r92JLQpNQQ3FMKGuDAxqcIKaz/t+PHt987
fTveSckLpDCRI7ZK7vrk9AMzSmQdZj/0yMHkd2tt8eUhQMNQXAqKjJNnr4e/J1+oYdY2lOSZaqBk
3idOwjFl5DOdrBo/IGrDrcav0jbkpkOjY+LQ/Kelc/C0T0m6P3dxgLlOTHlaStvwi/Emmm0FU3OV
nCoGvRJcprFTVgQ6Wz8XOd9NJRdXPRfiwt7Y0F4NItceskw2cqwzWALlUoeFqBbrQlilhthznQAL
UJn0rJdoVPAyezIvn3fKrlaKueCynPrBbLwIt6Afari8nKD8HySdNWnkDiTE4VLbR0rME2CYoIsm
oXR5rWX7RsroEpdT1nyk+/7fgAR9ib5JRsQVyGolMlBs2fN5kB80UcxsZXenF3dImVgr7ugtPbWe
Fx5dngbejzU4NipW9O4Z1HQbw46A06p3IFgcMap7Fh0RQzgx7tqz8aPjy4DroPFxbzQDs0aYABGX
IODhIoqoXCBBHt0hJsTXYJ2xbS2Zcet/P9H6xc7Y05OyPzSgBBYGLXwsNiTfIqYBmrNAtYi1GAVc
3YD8zZpx084CSUy0k4OhG3HwKstUY43WnMws3HSGaKBxVS5M7AkPb6UlctlC7e0xNsNlfUdzv+Np
9t3hHIUQtOOEZVRAsD+XQFmpekCj7u+luAeV2KNInxO8NvEAZs8h6tOrDVD0xoGqlzQcgIJJJWLA
37tH+OUvrpyR4G1SaBkHALD4zvebn8k5nHxEjhkRV/5slIDkoQcswC2bYAxrKQWxSip3jW7jx8sx
ee9Tre29DgesZrC3zdyVei5eapm33c9BYKGWyQ3Ha6DVjoJeEjjDPyn+NSBR7WsGnmtkxUZwS/z7
SZHIAJZV/CVM3XQcOGUv+KOFi5Pp6r3M7y6X5ipN5459BrxRoQeAu+DyJVgRMZMcTtZ4Zo10oFmm
uFQ5jOJrbVL4nuoECYMieHBOeI9dvQPk25DKNknSl/dT70nz0Hmpta6rjxR+iDnVlUT3t6C02bYD
oTxFf6mYeck3WTy0xfyERhth4sNVPc9FGr2Yd87SvSlPUhvQ6knLtKmIjYXP7VWZ8gWx3bAfFbaw
zl9fSgdkjnqT/eiy7ULImhQDeZ5eCnMtYhMC2jFt/P+JWxR7cqgM8AfXDW4DFZ8EzbG1pe9gx9Ni
YA8vHfJYEC4Q5rPkiUB4NE4dEnjNZbTJlG4+BwGu3OmYrlx+qWrdx9Usxzrk7lBfGiAXh6DcvY22
XzJAgU/XNBmiCuS18DzrEAbiirUmmpE8LyF9g6Qoq+GwNSiu05qSrjdj0kbO4oqjmcTBn00VcHck
aYIGSsrDwsybtqJrpDJs1fkXKGFmxmoJM7KaWYpboWK0nRN94aWhe9BjbkkQyqq1LYPfhPFVsBsi
Fg1+u8njUbqG6y4wqmuimVL0VdHCVx62TBvjDDYi4sH434G8xUrZHEBeOwvVGOm0tI6p7NPk3Bya
FMLCf/ftoOIl2C0qnlMaXrTQ96NrseIgugi6ypIRcbgQsCvvVOvOZEQRhwZWuED+Qg0H7MIPiV4o
fIQkxro6ury/dtb0yyay59ZE9/YRyMrlMr0aH0J1E1ZRlTDAIeGgJpnQ1bgC1Umi9/zuUmvguB2r
X/ngZBEGjrig4dr8wn98AzQCTV2AOb2iLwSZYfPoS0YmXEU8RupggsnjNGiVoONtdgCvDiYrtbDj
5Ssjca5l3oA0zLBChri8k/cUPHBzdKM9Eao68dIzCGck4tS30Dw8v2xUR4eZ1Wtr/F0ylReOpI+n
hWnu1TLLGqy1vanGoAGnxITFU8B+Cg3tfMBrBtZ64HninQu9BcJK4kygQm6k67UBAvhrQBMyYJYO
gGrWn/jt4t0XJf5ugrhMQ6Q70XR5m9j6Ru0XI2MOAXlJAwy1hzSxOO/CIIaej02RWsXYzhUfJTth
HsJDRN52Olva/9X57mwMzcn/7nITRGBxLPNN6j03PZQ7IfNeofNBizeDyvDYQO4WrtPSm+mnLUOI
hh1JT6ee8ENmhRCuOsZGdhVUJ80FGQwAjQQ/ELwBcrcy5OjkzSdDVmRa6PlFHmgYdk99y9HOxc4i
CQ5GTDSTDO79xfIjuqZYaTrz/KTRlfeumwB+LbWv3rDQ8VjWNDGuNFiWvFo63YgGeM0R495z9Gp+
eSXiJDIpvPe6XW57znRviylFVpBUFnwxhW2ImPWKjTZCIJOCRGo0ILI6ShrdQNJqIoEM3sh58q+C
l5p/EyWyZUW6FbPE3+V+zu9GJdaMSSkmT1A3OkdGfYi3KBt8skZ6CTvb7Eq9ehpqPKDWyxvb5Ur2
MrdZ+noTNHbZlsn7PGruA/E3CQo8Sst0F/1RYewY3HPmIsnrSRXG3VhsSTsTEH8kZxh8P8T3Rmve
jwpitweM/zugwu2Df/foXydYhF84xKPU9YYOKR57iGpuftPQcp3moCBnwB/nXjj3BlScul9sNUtQ
QzeRobHw8PBfPJiQeDwvtw0WiyzLsJNkd+26hjpwARBx4XLDL7oS0yOCGSKv6cngOsbxyoZTZUM/
r44t2rXMbaxlguIMQ7pF81zbCSYjy/WFBrnIzf4gTrUKE/LcXCVYv5SR4NjJ5xqyPeDi4+NqfSRu
vnPl1REAJWqxRQ61S+N+8CeQNOwx0pF/aBEqS809RF+Kbmd3W6aQ/+ArUB+zvx/MJF5Kl1jMlHn2
ek3rU6cCeDG17+e/qnUBkPgQDeo0PSw1rOm488zTeFmbOfRVAhimLH+DmgqOuIbtaR4GBgzh7qTz
UfOUcjz4x73TPHgI2x4JSBfzmlM6LHFHmxtil7Atnhi3dEqOYfzhMhmbWyLH3za+cr6VzVo2X4RH
y3MFI5pMGIa4zfuNLDBwD4jfojB93LJUEdKX6QKY+HoalKya4iAUQaEZXGClxg04Zhlgo+qWTE+E
/7PP6/rj2DMwmeH0voMj3EhgGBq2m19YHDaQTqvbSbzXBl0dbAYd35IhAUGUEILzdDZmQO7BVsP6
xzS4/oNJLzqW05iJ8QAX8rtzpSHx0qI2dfCO67GINMxuzueevYUbBwowG0pnqSPKRIfQ5L/B0Pyu
mrrxpvhENp4Z0IAQ6YE2TzBN4XiK2lK6JRj/E3UecDhPOHuayxpTMDUU7FICcjJPzsjmrE78+L5k
MGWbZyR3EUpykiZVvS1wr79iC3J5HUbbApLPM/ZNnm8U6X6Jm+e2ZsA0OjL+oav86IIDKGm8SLhh
7lB6/VgvL0IV+AT+lzlgu3GJ++F+M7a0gILQ1blRIlKKEDlsaFM3QA33QRcpxMWc/XjXIEhAYbDq
UAj6LbynHDMTkm3tngM7tmjEbHgzyzR1F8qFCw0K85XKSy1IFmf+Qsb67LSaeOjxiRUXRyFV0Dmf
U3Lo4topForG/ffrCG/gi/am4Ma1SxqIyM/RZicfCkxxV6gAAStasDbZOVYyBrAF6MZ+nV7AVXxA
FzNaLzjXsIYRaLH3QM1VHS3FJxBPHnDZSk7mahekCcmRga0/PaF+u+OXxpQmAGJs5F6gx1VSQ8sA
9FwSM2202Xem6Gmu8bdwHsBJI85cNP4PX81iIxzn+vFAGic1pzOUe5HBc3KG5Cs7lFlWq+PQyF3i
EwgR4+Yp+dZbXMIMZr2+a80FFQEs7KZJeApkvT/OvwUDGpR7s/zIjI6L+0j+j8+yzeuRk6MN20jA
tXMjPTpQKd6Sh/9lubajWjeRFsqfA+MhYPm3JUmdqpLRs/oriiMRHveHncm1hxCYmpoNURAE8DtA
MthYzjLZg+VLYKOVPqxIFyxaq5kP4ptjpWRi5/iSMfGjujKuKMHCqF2Q5FWp8aif1kT2Syh7xY1f
0VPwoSVAV++qZHpNOEEU+RnsNyw+Ord3/Hzfd8qEXr5aso4criyxFkGgzXREhr8ed+eYHAM7vvZe
63R/+wo3sliCJDYY6JJ/JSQNlKhNf5ndWXjCv7x/4j33SOyqSlm+RrWW2DCpnfk4caU0RFAKmboA
ppruMZ74zW2/rMWr1NaEcMbxsfJGKYhnP19b4KhG/Wuvz6DLRsH4UBquWDmTTLY2dfxV66k8VymP
sAmQnS1cHbHsvr2nG7/mSDIRUPvp5wh3VWDFS59cCc95Nrkq4iOxUnqJsHlHV0VEP6JeoBZ53Jei
5VcCO1hasrhLoLJo9BosWRIPvZcXk02XN/I5Isl0cZxlVHWNQlQl6gCvceJbBfphTN6uWgJx500V
dKIAukXbjje9Utd6Ju1vezcJ0AfYNCFIvRW5T1yNlt1WxLHYd+wTH8FfkpSg9sMXHJVlv1OUUpyV
Ch7UjU8wF3SHrWFxQipI1wxjx+AsKl04AgDzkJlhf4mJ9+MAsu/Vl2+FWvFJqYLMKoc+ViZMcRUG
QQBJPQFWm5p1UYwW/bvyBTf2xWdKMhAf7UCWOiO3dHieLYzkrbe5BB8gUE/TqEbQ/p/gmptbCzdY
qFnCevkVTsIXcvkita1k9psUbkOw2szUyKzv4Nf1W8gS2P25bGZO6vG1rxb+vVqp1KPaKgBI1ms1
DZhJlgJYNnQJboHbA51baX5WqODg4bgIhKmDrMFc2uEdX+RrldbuhRKGpHGTXo+idULDegEHiAJA
T21r9XlFsiicVmexGSEPEEwyv1t0izJpkq5RCvPNN4luR+peNquB37vs4aKgULTxrGmoj8qaNIIv
9g+hAuerMDWNJVFiF+GJCMTlBzPGPmDB09Uhya15udyp3woLFDf98r7p2S72dZXkXrDenSreV4Na
4zAmi5AJCxuCtk44owqa3+Y8JmFkFbDdNwdCXGLTo8ZU2sX5tAUN4rqeqJn6LKc6QM5jadPNKyk0
vymwy/0whr+yxK3YGEwAhJvMc+W9khcuwxaQXvi/GNQtDL3l66KB9qaqTp2G4TTvY072uSf+h/hd
zqDYRVD/e0EFA54OCwjf16qxbpvLubLcaAx0VgKJtf7ZL1zSTuY6OXMTvgfOJIIXGOLnDwsAORa+
50GBdt+XiP/pvyjpg3RPMWtXGsw41VMuDi4yVluEeakCGTNMBS9A3LZ4QaoGXBxJEC+9wWj6gkSK
arvy/3ymTxK4WbGtsNjZMNqXF20DY/YJU/OwVpKTQVTyirHd7Om0xJES9DT13NOqlbtnAKw87o8r
OzIdNBgLEfiTZfIZp95iGKR0r12K7gyInhhwste1/WT30cVivRfTWe9M2oqPrBObzVbqVtcyEIGj
o+YtcLaC8Ff7FvwdfCucVwZChTZAPlZhoPdwgsBHxkh0Lnnb+S0J6P3lFDQ0xh35bUN9aJd2o3nj
5qZTZxD3zZ4dABYjIUEaxayxabLgLgW0t/Bbspt0aTtkFxRntE3SUJHecCffO+BGBwZ/B6eCpB1/
HKlfa4o+KB/75WWOI8y29FgfVm+zyhEthbN0SCqBD2kQrg59G0Gm6QpUuFDa1bKBL607sZ86PKYl
m7GgqhcR3uZbuqj6JtaK2Rgvl9Ms6NDORhn7jcQjrBAbACF6x0n5OZ7LFO6UPb5Ux1ze9nDEiE5q
UDX2LzvUBl4ku9ao7KFwTUPvJeEinOEq/DKnjolZI3UMxigtfvyqoXsZBFBF7QR61k86pjkyCuD3
QYv3U/Lf9df2EKxSfi2yD01sjy79xol7UkIIyuV5QzauUG/rY3vZWDTVmqDzyWDoJvl5hDFds4uM
yXew+xMAuSKFpj+6qGICPnG5gl7PhFtR1cZXxGkrs6xdhSiFNpIZFlkg7T4apiKR3vhN7/Sxlmuu
0QP4fg+YgPp9Xl78B0Y8jx8AdfkDkiWW+Blrx8h5KAfoBIag6Vk5oUec0tZVPKFNm6IEn1QpbL77
5zUe5IhzhiEM4NC0nqZXV6RGqY72YfU8mFjDhTV6tPjbORrvHHn2TB2cksx7mN82+9KCT21EFQaG
9zIeohJEw79SM9cQ+PFsLzhbI0bzD1jPcptJyO9o0miJqSs36Yo6xX6yrBQ4G/tJw3oD+iRhrepl
QGmnuGvVa3n+2+5yipO2NDhR2YF7BrXm7wv5EcgRf5zcjjeTcyWbtBxkc/BWk74XJXX6wsw+enKX
AJYlitx362DBbyyUBiJR9Nx2WnsRPI1qvjx3TyeJs1dn5RscE488+MvsmJNjYlXueGR3wANknLha
JgAyBDp6DvHCc71VidBOTYBfmvmErC9ApmuxMoE7gz1QqaWgsgmQ2bJraXCd2rjlGeRReQ4y/DvJ
0OLdTNSovASaZFziFmtay+j/UuYuamwgBXHuJzf0te8gQ4f+L2Nx6b/hnXAXY5fJdLqslk5edE43
Qftm57ZX05CSY0JBh41ACcTimi4EnK1TqM0TCJ4bCxk2Ay2nJeb24rhFrFXzv/KYg56C2wzqnUNq
ThYyrOi/kjli+MBXVjsfbGTvpv9UXn1L24tLTBWeL1+Tfw1cXETFli7NIsQXsMT5mPhg6KcfgBnT
9g0oSa9nXfaI/VTbYSxpccIZKygTaFei2fMX2q11q3HSVd19t0/MA9qEd4a1LfbKoVHw0g5s8O9k
q44P0NsDaqwfiAalRg0RLgJLDVtAKlxXJQ/VpG/HL20ZZx+GjfpyCL/wexd+7zY1mnHgQJuc5l9w
j6CZY4H8+cCefoFmyL6KiLRODWU4chilFWCAv0QKNWvUTudhYvCJNglteyt3i6l5MKgdXh0e4EZ0
foZ7vAccMU87QgdBX1jT8Eox1K0s6lOAsGA2LOmmAgYqisxyWYzNYJzbwjixK/dpaGrCu9tVmi1F
3SKEOeI6eJTG2x4eKOMHe3XiMhpu65DL/AegARSvxbBCKFmWD2or1cFHABzHQv8aSTb+FwKw6lej
gtQKASMT6dQFknkEuRyhEPHu9/VCU4rp0AZ3auN9S0pH4YOr8nKaubePKt749YdPzdh7+B70w4ot
d3wLedCd3jdoeJTOU64vhOv2LXFbceFaLMpFlfRM40BCTV0tXaCrdaYaTHdB5mM942AetTzudz1f
L+EaQwQHqCrJTqBx6B74hO2FbRytNo/jNgASm7Bw1/JgEy8rynjWrfX2sIqLeipZNf15I/C4G3rk
+LtZGf8Jbgn9t49NoeSeiF1DUWIkeHli7n8Dt4Hxaw1lVccDvSl4FXslEOUrhJkSqciYBupI0fEb
EDPSCyPWTesZGAaTOatyEGNax6J4byW3+69+TeRLNh3FqghqYQvsfkWyMt1xf8j/U1cofZRj/Oga
R1jBsw01ArlGDhqPjq9UVgMQycCG5UISObgU3t4npAfsehCm7kAnr8K/zuEip9Cf+QIKcijmb8MB
8iOvzlbBfp06h7jj3UzHiC11j7erUzxLrskoQMLc6A2jaHBHIRjTU6S3m27Pu9EfNU71w+MnuOVy
gQ3YZeFAZS4jr9bad+9lxWgHCO5S5FS3vyVgwUhALMu5I78rs0OrZ7OlQjxnMcDG/0svi5/np2P5
g2J1nUnnzNUmAC0bIYaqtQ/cO+YbzDDksTSBx2u5amINbBICr6YGUyav+h+464o+Mr71UkFA+mDP
FyD9Wqx5c9UoOSRODPYHgZ+rkXVHoOiLHywuuhgFPICJ4w81AyQcbR828THQWPRq9wyX2N8Jyqx+
xE4W+U5F16R+SDixyU4b/52XKZWBPNEjU3lSbsRqz6B8gRc4smOmFtW/yiirPB8SnXmUXObg7jx7
2hui8FeSkY+A9ixq1SHEAN7dsQT8rtOh/z9bGcTG/revF/iD7KfNrlz/5/parLPxEmda6/PCjN0k
NLtmcEubNpLEdXng+AodskwK7er40g7BEvgsy6TLEC3E21HUyYx8mYy88gkZBTywqWi6pSuqcmsX
/7CjBzQSTXs8xEM48q0Y2nMg/TG4vlVxYctEehOTcHXoITJ6qPBjGi3veMV22BPGO9p8FBrSVuRa
+KQmYIT62zYux0Oc9IPD5LbvIXTRV2I1aQawK5PKfp3sZlo5Y84u8mNvJFoPTZsTN+7f62YcSLue
8oCXYuMaeTWUefz9TsBGSBm/aKJYewm9BfGSGAjSZNoyQowru2uNgCG0oqXjIXRaCWmEzw/78fMx
yefKzlFSsMuR4RY74ABFE6Z3TGqse0pBg3DpBE9vD1g5G4Zz1RQFPhl7ibYch+TQq8bzh0MyHH6H
BtC9HVY8IXowai7eK3RYJgBdHulpTUefEcPgcgOUHQtsfqcEkn3MbDCXB+ph0f592dty+yplX25X
PJziEovABY1tSfO/nRDxOsrFhLOxcquZofbEMQreYoC3A31F0wE99E5vs+oXo0kON9qff962RBA9
G4NqpoM0fPAxQDrO5KDXWfY51ut8zUtAHbBKyhYiTxuT4DoFUWF1Uve5wIuiYw2LXiHd2/Bq1/o7
xCMOLthjmR4gYAmdXvR4OEMfFJUQcIxPdstBNjO2NhYs8uVX8/ZIDJ7dnqEsUsnaBD/q8h0ypCYa
/BiCjgrjx4xPu/RaRwzUE0zcu/+hLvnHavVLCER91n0oc/7DpbwK4f5l5syTOlYxK+qO4c/aOW7v
w6caIZZIjuy54b+QNG3rhZN9ALav85ZaJbHcSqQ5oBSuQ9SUzprnq2xdF629P0f2VZCNR4WtNJ4W
cvWjK8EeFFzKjQ5lyFMTIOzAlKI/03hysskwn/3ryEDl4/UYdn1Oasy5xfLCzsu7NXPydK/qE/ML
ihG396Te+xnD4BgIcP4trhhsFaV7f806x3bghP8LgPKj+k243ju0XZy2UYfq1YOr6c85s71k0uJE
mQRyF7jIHr9yac5mL+J0Cd/huNemY6GCQi8JPZlUmvAP18rHloX12IVNfayxmmgrtIz8cZHjI1/Z
rblwrcuhKpv1MMKwslDukcLUGkZ2mI16Fmqjy+suU3h6puPylUXa+und7dGCWl5Hawd4rzFXrqvU
BFee0/3yJScsvr9w+VPm+1gJhP1H96PXdcHbWTkYWdWBlIMmC2sQ0BgEu+7uSkXDDip+1NJMYH/N
WSPZQ0EKS+SFPyqjPirQDE7uPEvDieZncCgLFUleDZfIBJUN74/IQCNtCf4GuIcoo8VybjwtH3Cd
+bzWbmiH1OofzQlaux2P2w74P3AvoY9V9r01nw4J0RIxHcPF1vf/E6P+LpcixDUZTxCdH6P+B6jZ
+VBLllkL70I2TE0mX1SVYqi6gnPUPsyPwO92WjzAkv7QBbDN33LyrVdZV+BMDXKX2hgNbrNx6vkQ
lwbikr/6anedhNlySiTnWtNbGJsiTVcSLq/wH79LYkZwcHUIow8tMO2d1y2/MYRc9+covpcLnJtV
BzPErgkgsEF2+aH9xb3kD8m9G3IJ0vVka8BUH+Q+CZVES8seZJrDezIY7u93IN8VRA836KxTgMAD
QbhYysBfQYd+htbEGexdLU9dpznTHga7TbGzgksLneZCkiHlAijQBHZpFYUQmbA+MyUXK1J0CUHW
FTJ+Cbq4cWvABQfZ6CMqHF5RaFWYjEeAcHL4ed47GhYYmXe4hd+cgptIdk5n3h49Ryvzfapj/zDo
e1YNHLdphaEhfkgqmeF51MEAQCUJxTbsjE2Fo6dzZ150ZZ9j/uFWMIjR+jOuCJioMajTpN2fibHU
q+yRsAfr14rCbSktQZfgX45l/37M9uDkQPXXoEdwMUcTK4hjIYs68/85+41q06bvAgKC0pnn3Qbd
NAPJ3WrjG5gyrFRsccozCDeHL8oEQz3FNwzepcANtwCF7qSNP+DvP0FsEk2mPB8lgJ7u0Yi5XXiB
oi8YL2xjeJUMshuSiRabh43luOjXFrLwh6ghJYoaJzzXUd3ksXuWCIgohfLwiQ+ygloVBQ+8idFo
uv8fL4XW4y28UYmWM2k/kPY4ELhZRKnNrW6vXmSeocLADETYawEMRhgIQ1ESwVSFJExT+J6bvAzI
qsZi0LXegLMyrfYwFyifcPr2njmrTMk8jmTpibxn9/0E0V89AyG6SKLW60kGvNCTS7/vz0YtMyCv
y4gXfFmyKh88KNoW4jiThuAPXQhIztiGAVz5RvUNWBy2Kk+p7wqrJR1P62vo/7+5q+G1vcdsCufH
a4PWtCgQuSfGf9H32iu0+rFhldTR9SjOtKNuHShqT8nY+FqQRFVjjWyjul4cs2bKCfNr8LgKEWww
Wk+ihIPDX1X8g2wVJuMhNoSFmL79BuL911q+tn2MlgqHr9AtnBQQB6QHGU8fmB1f8feSUU9KxHBC
SU93wVITgWUbRNRM5uROZymUYWt9rqeIyuo68oJzcH+YshBqcXbxTR7KY7DdemFcAOC62v+t8z6V
m8VGrilf/VzYS70YFH9+LnIWZuaNt0PER3+JnE7v3uwnhNvyBv4MiPkz4YMRNQ73AO/2CNKUiMFn
S9eaK7NWds0QyIQc3/ezb4mNR1ofPIlvFwSqdVGGILu9CegM9aCdJlFpCQs3EiLAZTEa8hJ8akUK
LsAVKmb18SduMJ9NadalX3d5Afap8AUThperhJaJM5HhikOsXPlWJP42coktJ+jPgkXvhUcgbpXN
Biuz7aOrWee9AotrP8BNc/lq3oKVPdbaUz7XJ6XA4gHcAzv5ueJEk5bXRl8OoFpVq7/OAjbZWA8/
nbNBwCqSfp3HFiYqmyZ1EOW5xQwj6MOMYn0JPOv9art+ZdJvT4//p7YIJqgLircqJ02sOTQ7CDdf
sLu2zp7hiKcI/GlHLcg1S+Pq9w1y2HjEEFlCuEqgMK0vZqfhtNfeeBFupR8XpYkduEs5gBrOKe8H
XPd5SqeYciMFfmKkBLzsYEFolP/h6in94fq7tWr0e7PmrbXStnnUsxv8Up0lp4OgiSfACLKMyzlr
td42F4HOppmt/uVzI+TlIULIXi1fOXD6R1oM529+SKK/oTGfy1FTPEoutKGADVmtwdf0MPt0ztau
AzgbO19m+cxktwYTTRAQXr3J04IZrER6C2ZzNFguYXGAqNzQGK8c3OFvErBKKrcBFDN52CBxvY43
bCLnhLTKCjRTpgWNc9FbqmyJGEZerjjBp/mujr3plploQs6iCkHS74a1hj1sn3E/3TPmVPX85Wvm
fXZt7g1ZfUzoNbqhBXHBmUTPjQfg6zf0RNWB+mw8gzvMzfaa20VL/Kl7/yjOpaTMiREJnphHr3CR
hcWiIa2bAAezERtqDa/cqD04zcEhdIzeqxazXzWtmcoutDSJqBPPV4IGvBo7cwSR8Q2nCLJ8hIDP
zj1KicHp0YotBH+wVDMiMZ8N3x9yCIkZtSjnia63BtFKUoDZHZK1QO0TFmI4XOymVicxEc2yuX4P
XnyW3Meo0ARuEoaTHqkoudIh0YHFaKfLw/qNaj0uutwOVnc8m7k1hFjsWAwyJEMbjlrxZAaWHSP0
/fTd7Y0JPRvVvm6oXilxPjgU7d2MGCq0P1V0D+1G3m4xMeBRxm0bLxJYkcvt+5+wW2KSK8cI1JNx
u5rcMAFL3/AChjGJs5Bfi7byTdiInUWTdBSw4j7xwQmkOswZbdyF1HYhwBQ4fNl84fJiqEp+i+dd
lglQKAjQ9ZUTqcXe15uxPBLYA/c115UzH8YJkOmvW74w/bqTMqhUfaA9/+IVByUwzHyuOOdkjNI7
huhVClFLlprA3BVyb+/fD2OKZgvM4tSMU9YJH0Aa4huR8JTMeZ+kBp5vfvwd8QFwejNBTsNMizuJ
szjLszoJlM1fZDUCCy4XNLFg37ROhUeTSHAO/ACkDJRB49XmC8DF0YxUuvHRH0nDNhqX1+UzuudH
f/frLYHCK4KMX+NZzYpDcpHFNt5WdmS9ZWeUvjDPsFt5JotKpdvY3RscjavgIa/6cmc1H0mDvWRm
W1vK715K5DFodD3/DuG/UEPSQNM8uq7W5HFwWhhMo2Cje/xPjwVQ2luwnShaCYfq6oNJtDLRVjjM
iiyuouERJvtgg1gqAbhN/Rrr6i06hOHKcL9jqnhpLs5B9q8aK6HBQV/UaMt+ih0DCnjHRpcs6Hay
lbqFLPqQUAdqCOe8BdCwXG3OPzhW87tWGdj/vVaukeraIlbOC7UdXQLvpIsUzvA0Hl0SAC/BD/CJ
iAmufGNUQUtfs1H4JtN6NSwDR+mTiuNox60lYydFUjU+htvLhKwbsSR0GrbRGRF9qa10hVy3QJTD
fItJf/Mg1aFiMNOfKaJZLMfKUBwOg9ko//Nn0HPdRPws4ScNdFsfe1tYyVOeXXpWylrZUFVysd1M
6IQkMSVIiH+J9q1QlIY5iv18NDTWVwciOXM+xW0JjjGzY6Ve8JGonUe6ep2qSA6P8QUilANAIUeJ
A8rFhnLDgvMLOFaijVyiUTAdPGeade5gtv1BnV+idqpvWqZqxHbof708Au2FWIZXez35ZUYOVY6Z
JfUvwCVtoM+Y9WQe9ZsxbNGyaFMBHLYck+6+4w7NDoNOxj+y4Vq1YJJg8Vsyihw1gFTCEuEwuUj4
1798DBtVqumyYaiW9WJOM+ZE1b0njemiycaE5KNgPt6OWGzuk9XOKEoCZHoV5SB3IH0Q/0w5cTZP
9uxRrc7IMrNm1uWbcwQ38Pl2LDO44bzxMW5pzAIliI5cPxTiiGZXYbvzW6KvT8yuBcXvIj6nEW0v
3eTDhwuIBAugdfXrGZSKhNHALtG7w7Tzfx03wN7az9JtEAzxthj+n97KJKnG+pImjM5YvBXPq7Fn
RvlB8xvWo9FUDOonBYinbFKTpCZ91FC3fE4OlYlFcKH1pQDewKcGV09Qj5Xko2dWEb0HwhL7L55Y
GkaW8BE9Fcqn0M49PlrU5VVUj94aEH2P1m+DiyiTLT5McWfIGNtdBa+kl8aqwnCD5NGetNz6eDYj
6yRxonTVgCYY5v43qtNtags5Yk+SRoxI+NYMQRcIrLzwex2Wgnbcxp08Kyt0UUf0kEXAntuxaMdf
npfFl9+Z1RjMrYuA8nnc4n09KyPeBDBgUDatl+tCZ0klSY8R6l2ztvQaBQAxmFpsp1XWBd91m9cM
evUw/4f+u40QKmTbMnZyRR6cnYa0lYmFEuFFcHLL66VCmLhsQernD8VR/Jl86NuW+lbwYltzz7ci
btNpB/2cou++oKww1fCR/DLmYMMHXN+3QiH27nD7T+UNimC9k2QVl/9gqHijS3CPtS6CNa3aVkG4
LRi/tZXj5TwykQPS85WO/plfSkK/JzlBNHIt4K9Bt0ynzUrBjaX4ztttu6ffZj7F653rWkTum7Ol
HCZkgC8tRyiDV9tu5JqqQzV7exCW99wjTHEoS7gEzplCK50dKpyNC4LQUBpbES9yU2woE7/EPptL
JJSo6aPfMqmO1HFIX3L7iKvMPARPMM8xFuXk7JQmda7uzV5zj8nxycUvCoLWARsz5AFEfh0cHy9q
aZXfZ78TCFtYCvYZiIvVxnbFu5WiaZkU6kgZAnVC+s80TQMlvnYNMqrwKcARXAQVhUh5gIaO42cW
Pm7pX7Zwfr5IRZqMnOmkYo/ZwENhN3c59w1IdarmPPyzmQFMJ3upT5XO5WqfNu3gAt2FqIW0qXsD
DxocKyh9YBMuXFuVDx5NKEFogOJlQ+H6gX1BBMIfxvO4dOZMAwx4sjM9qZTJK5jYoqMMfqVZXrl0
kNGIPxSQypeEMnaKbS+OHwJ6UsQQOf3hRkDX3l3LKJPHrWo89UDubOABfoR71vPGyUvGFPj/FtMo
Zvi3GWGQH2eVr9UKN5xkTN2Q8ZoVdvZqWFgQvPtz8qy321nxaacXlMkdFKZYBfu/dRWlzUtifIx1
h5/P6TK8K8ihSx0RUtP9Bidcyx9ovJQwBtzCMentT2a+rQvXFgp+tZmW9UdkVd6TogohR56x0Zat
gvb3pxbOUQgiSvsp+TlBE+IYgM6ciov5Jlku85XnUJGtSJ2e2WQYwiYpK7cZd+Oydinb6CwX7ySn
aw8YfuMV336kgB50vJ7mxv+h8FW7dhSJlxa5PpBYax6ZHQ7hYYDsJs9b6hp/h+8DjlMP1gJdLBVw
kYoMQ/e/IH1Ovg8MiLDVhUe7wrrv7WpS8fx6rGg0P9zNjgTJz1Hl1KXXO9bY34FAKuuMxLu7q8K/
7vthjsK4lDNC+xVcTDQFvqzevhv/2SJwB2jHuM8wrLbDnhk7HNnLGGOnbxgXchpIZGPZfJFPwLQ/
mEHf3do2PVPvJTZMAOKIsQN1xBF5JI0zrKJxxIojwUb5x3zB7IUAucClKK32uiB8CQeuofdIbXnI
i+DAfPbvNFWPzhLRmRagVb1RVFmyuhug/EbaWlwMB/sP4p2HdRQYKO9Mk7UVUZbKy5sktR9DxAd8
LHquG6e0RiPe7qm8qwYEizh1pGJulRwS7Xdgxnl/+drxRPPkvgHaQCxtkSu8EpJFHUAzzdkAeN3c
js4Yjeugk0r6IJHniQVwfSK5AQ1815Zvgw31ss2W6tp1rYq3xnKurqEoeYQOoOZ/X9xwlIUisZBH
XwNKndVlQtLhXd4739ehcN6SEs/YoPN+IXhiii9VjIPt7C0kh+itRjujUNXcrF3bzIxvB+hXcSeu
YmFhBIODQZjZbMpMBjjor8UjPr3HNIaB95SOWmnOL2GyRYaMmjdLvsnh5LSMnsCZ5YKbNRC8g4qd
0fHOrB/GlM5G5DOqosCmvRViHAfTtuq+TElZDxZnKrIGYwFa/P7duLfN62S6cxgtt1NvzgjIVhpa
bKBOLQBKjzcfHvP9xrwvkPFo6NeBbbj+pq0SapOT0S3tSCCTNkIuB0Wmtb0QZvjvgNaMqTfFwhYe
BpMeAYPMoADFAcUhA4VtytjCwgQO3mQr+ePseiz0PM2Ct8EkQADS+hTDIRtta5nBTpqeSc5bswmf
syIzUUHje30g5NVK99w30y1Gx/Pv+X1acU20N4ykRYJPUxlVXVV39fdHU9r43WCorju6taPyB97p
o6QdJEL5WQVgmQS7OIRclXL+pMFO/689hNf1WagwQS4MyDjk0DRwrTgRxUmoGtSRJ2RiQdfxoHf2
tsLI3eZQ/YmIZvHje13WTd/E0ZGsnGHsbKIBr+UJT4GZOA+X00xPWrcn7xrUXNBGVWphXZ0Y82SZ
Fcb6NsLmWaPpaeuABXXwAWMcc/IEt7PnVbiJbOaGhPNMoToUjxXiK/EyjDTBQSXke5jJgie9EDQA
E8pc2RW2FSkqMwtb0GsOwelouvYwyX8qebQytFNRNyAprGitW1LbdFm1lg14jhIqFasIdpZXALQG
34lXWTS3tS1dUzxaQvqbWaueXyxQXxhobHdTIubtjx6EJiIWvvh11T5lTPakIikxJL6KMK35cWjV
cEnqJfsKAX7qzva9TMZvLsm4x6F/EtculYlSyhtJ2pHrDE8sR64x6a1EK2xqTgtMTSQchCNOu3n1
y7iZ/dTQ4Qu+N0S5mVnY8ioNMIlr+RmawWEBYXisqn7FrmyxPGLGfcii7JV8QkAJDZt6wWIRdDhV
z66qMFiv+av3bN61XWIqJOj82WWE8r+tL7PSHAkPf4FJ1pQjX72HgY5QjxkP7r6ANjTjPQEvM73U
6Au54erTruwKS6ir3qaFl+iF+tLY3opSq0Tp/TJflVZlzysSY/m9nlQEyIxcWFlZEH9+3Nj6B1xK
5beHmNT2tOnR0tccgX0vEo8rgu4c4cjkx6MlGornHNEMDx15uEky6s8OjaR8ju+NFGzdtwka6p7E
IHpH7UVTz3daLU9TmffcMrbO1z58xFqzYzN/pXRR1yLj9Xro1+pdsYvuJOHoeo3cpeplFA/fjcKl
UBtXNfp0iXsMT8VM0ovnDV9k+wHyi1de7W6UcOdfe/kqsuE8Mq77VcTxKG6TT2XKxdH18dcOXhH0
ZYysG1OUEGm6IP96G53exkZCFIvh7EygrV65xxM9ZIxnpxsFX+g5mHcPzGaD7OqQR0hHwfqeMBSU
wShtWDAbpk+gUFrXlOWKeV1AWfgo2DNEialXqYMcJkksjgE09a/jaXj+8kXDcGimBjzav3pjVoie
T84IYe7zAD5pp09BinbPKSrojWqSHTHeKu2RUVJvovBNadd11GStK0nbBmiY/QMccpzyr7SjoTqG
h4Vc+z6S+6v9BGrp447KNSOjPiI4042LtP2HTUYHmwHTP6HC4Dw1SbpIumlwRfcPg26x38C+G7pH
tkHtmttowSE8GdGVgvNigWc/3MQNTb1shz8RQEbPv8rm8oUeLvJIfMqusq+xsRJHDebG4pPOHlvO
7uPb4/Iv0Fzne6JQMNhXvtmPTvEc4oNcGGitMMSqSwpEBWSm9yqYh2/pDZd4fDhld+0MIFn8uXzc
vZisjxWC1BtEBJn+HmsnAoBdRISmREjPXfwMIwb6LFGkSYorWyY/rfBPBNUqfOcSL6uDqV6NeeAW
Pmi3MF1e72bts2L9kNgxw9xwwGIEMiCfAk3gVSU+5QPHQ5elSFY9M91xlfKUwuo6eW/f2Sc5Uc5S
gIuMm6lCeVTtH7qmLdOwNQquX623foIJliQ2bDwibxTwR6Pno2k71aDKwAicp8F1eSxGQ7kjyxkA
uCD54L1b7R+6RKy7FauHr4Htvha5Vs/0a3On6P1FppW6QNIViG+a22UQMvFZGEyWd5j4peUBRQSy
q8ISQL9Xg6WnnaL9z59QUA0Uaz/6nYMfL+e57dPM9WsDQxrrxJl3gmwU6neJP/Lu+Twb4Wh1TlNQ
Sm1sYcNrinrLYSFLigbwj8q1JAUxI6bct5d47ScvheaKimN1eAN/1s+f5TEDM7SmTSphv38Sp2P8
k8ElfnKPBdLyGqhV0LCcpstfqIy5GIBIupaFx/WeO1dhnARaRFkLUgi0rCB3bLQ1nv5fENnWgc8R
PL/Y3dov5fvH16pb/pp90ZPHoRRYGlbf63TMTgKrr5tPevqB3b4fyF9MtspUHHphr1QOd1ovKt9v
9WfwWuDXYxUTeb3jILJKt9ynbsdloSEbL5yXRbkpEcKqNkxg3acEFZsJOycut2wFJwZVLjEpYZc9
8DWjdeUsKuA76ydFxVVNBisjd1ZLDix2rOFlsyAP7kJru8UeXGcGImz7RLAVJt4aauk/Ef3/QjJi
zmmV5oxqiJltKo47izN+WYeQtrMHZA+foWBZAMO3XIsuT70yFYCRiutP1Qs+bYRfjrP0vzNkc2wH
XBOJqzr9pSmPKipk4XFz/pPbr1ShNe6PDwFTosTnebjaZRfUQ+NqqjpnscKTm5/wa+Y9j0stisLW
Xkz31PUseH1FwUwYMjMEikXPtjfF8TPCVhMHEDxcWbpyFaB53YoDIRj2LcwUFFPUzHtpJtb0l8AA
UgoWQe8jzksK78lxR7Os6uyU3jE4nMTWRLBKSjd07KoYzyMuHiYHxa649JMDIb/tKRR8ePVs5GBw
vhomSjypb1q01Z075fagyBxWBaeO2uEnYrygVe0c1qd3Og4nSu5U2wkqX3+RNBpGYXBSlOWO4V6E
BJryPt3gVDjRexzn2kQsp3xBgRglrz6exdSs7Vor++0EWyO/OV2zWVz+1mXbTU9Vt6dstODWO9zV
1/eoJf9DBuUSSUUsgiyDafgEO/G9QhMzNFc0x7AzepBY7HsknQq/l7YiscjiUqMPbfOqI13I2+VW
cYuLW88dE11JYDjNEFMMGjbSmQF3BLeDJzwA1rbAzjOQoEF0eLNt7figf4XqHwngbJQqoxvBznVw
/Mkm8GhteLLPgFxTlmMCW5GuXlZN1LSf9/Hq85FnwqICw0AhoTvM9oNjMuYchgm1LznwnEVyfa8l
dB7NKPelqEoc5kKjeB3YdyQiOoszfSIp1535e2yEvv+DzOr/KMYrPRMkA/dcsxPLvlPFN1NXv0wr
gJaelLHc8Qr1suJCrWv0+QB+uuKWV1t63PLtaNWek4+M0E58j7Tbr+qlgzKYmfWmGoGxyAB1eQdq
uM1PmN5/ff7CxundK3GM32fvehkmkcpWNE4g6s7NKqhCsRIZbUwTVrRIceQ7F+5LC/0So2SvbVQ0
mHsf4t0jvzxM6Yy81rkj4YfaHLy+Typ3xvztet1tZtID1ikTpAWhM3NfkvDsLzL/F8M8THhVgK1m
LsQP71zhRADaKkq7ixi5hne35oFObtfqKQydmYYX4q+0xItvkbOEra03MTDsrTtNT1ihIbwWkwm+
qLJcxxWMdEJ90Ur+DRtZY2kK0UxNx4dPwZ30mi5b1Mcox9qqzECB1w7nISvLYKP1mMkWGXwid1CG
VtDKE06Ktw2VFwEDX9cEFyQUa0rSfhPegwiLRaSgAwyshCrPXn1NLnaRq6KSeKYz1mifCkpNmzb9
yby4e9atTQSNc1mmRqvBn/hOi6K6djIFDdF0jFrjSKB37C3mS87Bs/OAImR4eQ+JGe/UoGDY0Lpr
xDb1bMm5E4qb6CumAVq3J/orzL9CP7CST8/p7C4LFYoFlP5MLOcF/sZ/bl8ekSAiBU4X1CA/UhRt
PawBfTNqfJPQqYR6csHklanf6pPPgDZrwVOxhBYe9a0Bmeg6hkr87CK/R7i1AXFZ64KvFiQKayNs
bIHybDIYTejohZ1hEC8mylakopVBH3EzUZllQCYDSwwpJBMRB1E+OkcE0rz12cQQckzRTKN/RFEb
y3PtXk3snSTAB9ltbF2kr+sSl7UQa04NTMICpxK23h9czQUzi8RUL1vXH8y1ZHICwUA667uiWjgi
nbmoH81hV2pmb7Au9bthVDz/SLFXhy8v8/4AxT/R8AOs4UNAkr3E4dC6Utao8dPfVZU1u2y6/uld
G2t6Fz7m/IaqUEaV0M80DvL7yzTRNsNfJVxFsxTWn/4pqruoF3tLOV2WJSQ1y1z6py+fAg3aAS8M
VSH/dr6MRFHIhAoB2dEu31Hj0alv6tjp3rpQaswcJG/v8AfdOMVF6PjhfUkqns6DI09J3YUhmsj7
q+z/A/rDjKX8RnvKvisxlkFQk5QpPrG9OQPCIirWWmpjBQJ8j2eKAp4E2i9bxbIat/6Ml2d7TKh8
foQM805dV8+q+3TQFpplzmdlVABXbQ2IhDvAwIgzbK+hVE26EgTBJk9t5SCxbkPC19kF5uhFDPo8
EOdPghMnLVaJSO1k4W/Bjj6Uv2FeapiBe/qWxnjxfqpVXQ/bXMWaQ8FZZvDbtAIDhd7Pp1IbYv23
lvqGMLjdIcNP0LralFZ9XioDay6LC+bnBkbDsXzE339z3xLwLvQf2uh7734KC/0FCVYNGEvwB6G1
eebTfsVFnQMKoraZZTReEUY4FWcux4oy9n1F6jeJ44AxuP3umo9T7NglD7kIOXB44dJ4rHOp9sqw
P/vp5vAtVY+yinkx4sqiZiPPV2/fGPMgGUS5sjKsvwGljM6OGsk+5AAXbYD4NfO6NSZ0mlbZKFIZ
1kZLqcHkwZRTKhOdG1jF8jLdA6x9eJ02X5Mj6GU2KuEdi7vvqeGOYaTqHbWb0KciDwFPYFP+ZOnU
XmF3mCbvwABho9ebiViu49S0Nyx5UOkO4byuxDyBeS6A4RB5fU/9dIwPURHq8VFxm4673MJ6FQs1
rd4QN2j8Y6wlBG4FbCBn8paYdLqA33zXIlkoy1SxpasE7rN559Uqf+/XR5h0z3d4YjGoRj1QLC9O
MSWcFR9P5sqcIyRhAMy3lHzfar9mBYS3og4VTO2Z43LJ4/WodvfBSmghwOyOYUJy/gxFVIHkbixe
iBhME45L7FEmIlo3JkG82NXHhGYaC4qNHszXhrSyhe1dy5jbcTmZqNAiq7ddhI5Gkkyrx31ZKqHt
Fmji+CT5ylviKBxPB4uwLJg51G4qT45z8S/jwK6JFYDelsLfb22arQhlXlKzn86opBAwNSoek0JE
KsBHe3s75KdT9fTqoW6mBtsrvZyqlyGdlABXpT/wPWu/KMvCm0A8vQV7wh7O0vm/mMz3vVqti5Ic
LOb1aTCV2B8e4eyNkJ80SLcgFemWp/kaAa7N66DX9IF0eIf29QjW2y4TT9TeE/rGX76qTvASjNO2
Ukz84P/F5qHERw4NgKuqCC82sI5nsrokPLa9eAzL42cv3+OzIUR/7CJ4OLu8ycTB0d+mJGkpGezN
cVb/BUv1PliVqP1Rd7wjnFESfIAN7QzwI406CYR+rHEqMggNOMcJF2lwiyu8AZjK2pxRgQp+cjU2
D3+OFwEtkjP1BBF5tkaLDMCooDxuwSjTeioVIzGdpr8qYQN5vHRMuXG9iiKD/O52dmpdLgKPgxdH
z+ZTwvXEnpUEvyBXy8F0u5u75aLn+eiXuEoQ5p5W1/bqH85G1hjXAJGw/No71plcj6gzRKxnfTte
LDxyBwrNAD4rTTmNr8faU8+ojyCWDcUSKsnNINPn4hepw2rxLSuKKTt2QYM2WSidanAMuf5csOOQ
HgZ8enh1KrZxCqW93t8TyGmkZipoNFnQKFN/EhBgVMarjw+Itpacisk6desqmmvagm/IAAKxUNJQ
VGkJoKEHM7J3auxANDjqnSNSsls0R1yZDCJD26lvbCLetnjUNae+VwIlPb078WokeU4bq3TD1Hx8
I9f+YwYLS74HCvSVd4+JFkdKt/e+by6R0mhdE7tLKvMR2/FEzBPXR2cdJGTfOK2aAcRE8oQMrQwF
YcJZzbzZynE7O8qZhR1rcoSJilnpX1znFFED11JBFXaC29hXMkQBwnSgOEDQong3H5JGzFL2xsZE
OVDlvMkqkPsnlfFRP09BNep034gegILiEW8BtTicRreNZUH3g5dhkJlQk9jo/XREL125oIJjAwG/
N4UVCnJD2ot3VR06qlzXOgakgeonA4jbTFf3GuvcqB2cNVKkWwXwO0zYFCZ7PudU2/v/EP2VG4G5
3oX64EIfYECSaxyOdcoScvs+A5ZET9D/FzxjYn1vcujA7v7KzBBIzLlGcqXMqUNFgrNgjiJwOMzg
OVLUSsG3ldNyKzxuGgYyfwP6LgO/GXSoLXTYvVPWO6qJD9hSfeqBmev0EvFaVwP1SnDKHB1EDVaT
b1lUNXPf76vxJB6oKDuw6s1HUz8x9lW2ZKCR/oeyQGYatJBVdkViVfhXoCUAl4tLIDZZfF5FK8BD
dvLTAH82eWk4UvX2UU9M2ZGTRpBG1aYXDv4RZZ3OO2DCnA5glU104qyW9qFqWJBhxmaD80qCNIfA
xculTgiXHBgW4XLW9dby4EcWZiTzUQaEdRfAxFXXP0FM0y1VJAXXGSuXKrd8lXMQeLNkCW5cxB0n
Dl1ehmcGQrdi5UmRJG3SM/G9/ttRAxAtgQKKfxHDpWqKQMS79aAa5nVUeBGJ1iPYLpNOiJ0f6SEC
IJf6nxJQLF1TK9FwNerUd0TEKW+srfpMwYoxcCECWKWfOKKCwM3eR5aXRatH9XJKnVX3rrO+UL+4
8VhUst3t1WzSb04PUd2uPL7/axBn+YZZ4lQGAvkF55D1MJfIAKsu534osBC15SBGC3CXXlPn07lT
/R9eox3lXjFRPM7t/EhI+Lfitmjv3EpIuT5Tc/kc7QcDfBBJ3ehGJZ8bttP+Fle9VduVhMJbdohS
5xBF25zXBsNYYDfjZFf/4F7NT2x8YzImNc3PIrzWc9xh99UBP7zrgsnDqtrgqX26ZZYyRsUSAjV8
qoplJzoSgi/JuWlllKAqhOGIy3i9gjT0NSKLuZbChokz4Rsqtn02b9/XzOeB915evDoZ5t33WR1Y
hf6VKrNzW9WURC24pm9fJLakM0ddsO9i1W0Nj7zBNVL069og7PngaN6krwRQKzJVRZaXtCuO7ddO
WxfkIoqq/tDEpW1EFOxDnJPV71yr/sjRkRUP++xD90hQniy+BvOz0daz2xWuud3CxYy2w+/2Xcaw
kuEXtj0qrEQ+41rbW7K49tFEXeW1xPlqPhJJDQ4ZHMY2PZBcPC2YeuSZGo5u/P3X9yqQ2H/yGYZK
wuQfVM+CWgNxDyuH9VeHHTf3MtS0X4dW6xxoujK4kp+6wgyO8erH0GhB2PJfOvYQCBUup986jX8e
FelDfRAFP72vKchCRNWogT2SsS1MPU36LhW3BRumXRYUZBPgbXjNeh5Xx8ANIr4/rJutqWEGHd5c
0BiDS5ebSWqMO574F9h2JwQkWrMHtTYrQ/hUsvAnIWTpdyXVY5YG4oNZ86U5rgsl2TeH5AP6GRfB
ipk0Sn3hOnZjU49ImSgPZsioffVDborK0gzlhynwUAEbJRM9UTxbgOnRcZWrtzjePUxOQzEOWqh+
ksG4yv82FslQ6oXLTKWykjDQ+yUrYQJ7OlhjpOXiXvHlY2kc+m/lOdvp/lZA8nsDRlR2V44jRMtp
i214UtGikHF4EQxablDAL2dOpYBYvbrL/9VebYik7tfXpgD7UdbE+z8LwjOd5+V0omeer74o98W2
JwtTBR1nicOgpFKmV50szUPDanm1wzYW5jFjcFk/S6d5FoEi52Tl079DVMobUIAJ19YJkdcvKptv
4HcMhMT+ynCHo/r7Xc3IK6on32N7464wtlvjcCYELGrN+FQriv0gLtuZWKupNyT18HS6gWevKT2Z
7ACG0A2nq7akHrw8yVBPYPvNuZ6Q+LVRdRBUEHz65Ewnd4ADB5UXX38zbebUafRoCK7apGpuEDfL
qzO+bdnkVGUd8GOuvnNXdi4VU/7Irb66V81tId0YUuo9ttBYHeN9QqWxXz3AdCL2PXymoaENftMC
4crMNqgGTThniN68Aw+TFfYbWzE2FhXHahveufVAYv2SGmEHlCdweJ3UcQybnkMPfnQ8WhJA7SyF
0IkPUgvGuy6T93KQpM1xMDBnjvV+OJbzKlExuGt0epAqZpx2NLh42baPLXbu1CmYdFA6PHLPtRIK
4M/0CYYzEhOvPk8qKM7fvfaWlSNB2NyCd99zwcGUZUeMGpTckU36KYBXON62MMd3mEtqGNAbkSOy
gVRNFCflQabNTatTImuwKF9pktcGDQaxYN0EvJnCcv5MN6I0hqXphz+lBBOk6Z6s+LD87DC9F1c0
6FUsj5KKDoK2u4qaKskfTWmfQuXeu+qcB3pE/3q98+oqpOuDlVYAatT4wWrpOcjbDIK3jdpSv8mP
mvo/mm7/yHJJ4mJ5sKwnAgIcxX07J4r2xXTtdJ9iyayWe5lR8EVNgRKnIDpL87cshrPUv5D+JuZG
xLNGnX1YfgFp3eLvnCkJxarVxKrXoqldhQuKMZRdd8ywzp9IFdFYRMz3/M0evGOfvC9mJanOg4Q1
wOSuaPP+0otgBJQQOJRpZb/eA2/J2svdxFVr5MlCWGfQzUc4zxkRnAQu55KKEe5F+DLY1EmR2BUl
2t6PIppmp5ovr9XSJ0XEcxpOegS4Tl3RGMKSvAv3oaeGnu/V4wM1MhOzZ6MTLwfWf4DUERTZ9V/a
gyIbxkECyNeg8rLoiJDdyp8+AKhoXOEllsAp66GjeBfNl7qUlaA9F6b9yZLKqzaOQ9OMFX6ds+wJ
Frjw65zBYsq1rQ3Zo3HjRGvEONptDOikd18xmMasZB1cdprLqNW44auYZ8jpDHnnQonH8fJ1aHX1
NKQxTbXPwIqN5wTFhjeL3Vp5T1QUiepMxsJZpXlXtXpwazD8muZ90JNdpKC5HPYDyMxYJcyZEQXT
2pvyQJQc23MHjsAV1CczxpgxF0PD5RRH/uB1yq26Jh32AIuUADWIciFmKaBVS/mqLHEa5J/5x100
JmBd/U07TnlHw+JdLsZOeVEveJ/vH4hX5dVjxVnyNp2KKYLXjMN+5P1Mo676C+OcctYnxaV5eGrJ
V8uHhxymthKEOESQssNDXrAP4CrFhAs9cBsZmu3f+jT9FH6AtUf2kXQvh8PU6W7gaaB0GF6746Pr
9trQQ067IszFEGJcNMuVK+z7uNRJlWTs5Ssyyjv7KcWhQbq0naMDFLTCIxq1EFOXhmKdJEofvIbt
O8Ca16QSdDI56WQG+tDb8ehUHTl/GGCBFq7oa9UgIQNIkB4hQWyOobFGdjLCHvkmSV7hoPdWkSB/
L5H5pYZKfr68MdQMMTpr/Rltx6cnH1il4p9MbnDCAVv5+zoAksKo/u7kkTPiSFc80MAHeCIPegLd
B1AMdCnHHleg1wgaDZB/QvRn1bWZig4iuElrLZUcxulV8aKBSm0pPoQv8eA1ehKgF86WN6j1ioqZ
MbCu8iSdLhAmugR0/V1iatQr71uIB0pMggqIbxYij+kGfXn/JqJGS2xlHr0kXZIE5dNihkeTGojk
1gAUyhae9Modp3kOswTXiTyxToE+wgu4OaDLSXrCAmh9FmerVFWrsS41KAl/ZaujMSH2HgV/e8V8
dY5B1tRAwxh76YfpKC8mLd2AZBkZwBkljTmpEP2Wg1lBg5Ff3ZAwlO87/hsmnX9WO0t4jaIE5R+V
K4foJOena1KDBLGaoiZq443BPxPqQxiDlZ7BS/XcvniPs2pVsOTZf87Fyf9o9bG1+p9gdIU8SqW4
1UMlpM0c+yTb8O1iNAli1hX99+IdK5ws/xk/09vdK5wnx7Fcnfpwx1YkC61dZKkUSmWbxNQTRYX5
OBoEg59ICDBewjKQqx3HN7qsdCo0SI4pKxvv0HuVmC85fEVZTF/EKUajWEjMYB8rkFvvavQLhmb0
7ga6JBcMR1YXq1Ho81+Ggsom8YCPvUS9AVpCQiGDPY3CVodV9MCWKduohgdywn7pfQ4S5D8yrTW8
LfJuigDSn+cczF5SBDDEH54NnBl+/PDFqF/FPQ78DDByyWhmyMUdK02kRB/g7EBfIsR4CKIVNncH
Mbn7QbrxrudupvRkL2mV2zaXvkfvO8N5UP9Dnt1AZl34vJ6I0+si3CDSIywm/XLgLXTIZQWBhKZG
RhNPkU1Y0h3pYN8z1s9RsuhGNQ0oxJz2o0Yrutrz7eip+emN0klfwG7kEwcWe7AFTWeQaxX6NiU3
TFU2Z+p6+5HF3wWUqyox9xi0WH8zLqAmsxLvh/y+q5iAaufOtCoYyxFVhEvC3kow/KDg0wa8oNeP
AEyu3/qpOJ+NmBWSmHbC3E5Wf1J07aMuVM6rdNErITCkDxbynbGNycUQnHOCM+b0QqVPL6QbOPdc
FNG1f+XIobxwUTg6wwibWpnwV4aIL9Qjvua0XkltcgL0jZoCX3uK3xHrg1cqKw/jYeZCDyaIDxue
9o4IVMRB1MHRAqowHKz/LEFAoIfSbTagggN81M3IILfPo4gtm/GHbTDBVU9URfvNci/wDeQfTJ5i
KYx6YMiUZfhRlI7g1FLTveflpwdeRcKu5Pd1cWYhHGMHcFK6dxsj4FwQ1tiCSGdH47bFoxnaq1bC
JtwVcjQvinrWZ8oLOg3irpLVrxPQLEQy1RWcPNYr+dYP1tArrmJEutva1XiPupRpl3oQhugy+c1p
HwpNCl2W6Dpx+4Dhjg7k/mIWTM2o6rMMTG6EMcU3RG3g8wSCMhim/C1RmfpHL3A1iDhSWgi5XhTa
zcNwpr2/VDGxLJsUAvbemgoNR6yKtPtl76stYdjnnvxZnkjaOlHzKtP6pxq1L9UjKERnmKf/Fo5a
NIEhdqwVvduEFFG1qAU7qJgumwZjToaRG3S6X9OP//RJPYy9fUmCjr4R/U2a89ppJzI9+WV+6+nW
XsvnFnkEcRo1Xy7+6H1bLd8Q00jux3GagHdihS0A6Q35cU+Kj1GFLEr4nf4loWXaDTWuouaPDcaU
TVlscsBtKQIwKE2+h0QRu4IdLkuEDcDpVQP2ru3t8LanCSupVEAB0c4An96F8GXBJhaXXUtcwP91
cfZhs/H0NYo5TA/oyW5WDS8lbv6yRJAwv1Rzk3zs97ll3EyxDdlnXiidX5axbKEHkIRB8tniRFOF
pXUjsDwCSnGEL2C3U4HkV9cFkdNYv+tk0t26ugtDDZ5m156E38JHPdxTLcwCxktLlAQyJRFDVQYn
NOItQJtd23I2ErDNmMMB05OudCQ7F2kZzlX0sRtCLA4Qnsdw7OseZUQ9sg6ABrDfQDDBRor3Az/9
A4cH5+6EdvIBF/V/KbxYpo7kNUljOEzDaH1xPags7VDinDETareT1akrZzqTg7dwTZW4mJ5JiaRG
hps2+EIQADKcnch//96axgK9fdlmRYHBKEA8ovtTnIvrQTwkSll57BVKgYlZM9pZdxYVP1QDr3j/
RHFgFY0aLl8cgMbmiXhosUO8W5DfbzZzRAMDbWKUgFE28jUex+U5mlE0GZXcA0A11DXCcoTdkKGA
CPt+z4g/lJogkRtSVYWG1m6jDG9saGYER0ay+S1zzFkqxTQNxEMTrYT8gOfZOscjc5z0ni+/UP03
dL9LEfNvqIfZz1VwNzfWytXeVRFSRUgmyk5GqoIZIRjrk1/k6vu8RFXdCs/0ysyCIad24fZw+XcQ
z3ds7To2EoMgP4m5UXH74DjE/fgiROAZBInIjZkUnPLaTftD1FIPK9RxU4YP2IzHBuWVQIQl3Q9A
L7x0bVrjui3HqcsJlJO8LghrB2Z1S0kQtTK6RzvCLVGE4uMLqtKK/93EckAm7XoQQfSaxtGUeqrO
armx4xQjmLoRKRjQMf1yfMDNrGwWHJtYHKCv/qwLVbx01Fi2EysBmB8Ctms7sKFbczFUJyRbyG20
PthrROh03uh2d5a0H130OE28+h1YLOr8FbUsZTfKXDtwodpm/GvluTzlByapryC02N5LNFiLJ9kY
3k5lMO3KdAlkrUhK+S8AXINBpSIUTGgn+I3mlCpt8X3aKogum0i3n2U169PyIdOaSikZbzFhIRnI
9LCOyERrNiK2roa0aCi4rxlughrijw4CavVQX/PHsZeMeHUbLpxgF19uTpIewYC7is0SAcXLGQ8k
/RlbHlYpDAGvaH8+MEnv2rqF25TYj8HynK5Mgper5mHrvbzj47gU0CQkd+YejHYyOcLhhHx66eCy
qs27UpezuU5JKvsgVEgjGMwXlEiGfBBM270agkWebpzaF9Gt9tytkJmJTyPsApdzhEKCURvuXC28
mwp1IHuhOQfTMbRdiOnGZWigHaKtLaOP5hHc24JiIpuuGdODQLbFDJRLFq4aRD9/SY6/4fOu0Fwl
8wkaHh6Z1lfPPPW4q8WIrijLmPma37ql8TyQBJzI0wq4MKkF42wHYNpYaSU3R2eThjqrV5jlvVkt
0kEniayk2yGoFSdtaOzEznmIJrX7yJmw4ctGDe2Q8j/9wBqeiOIfXJawq/yBXklWBaxkWI3RJ654
RD44PmgBCR6Gi5FHF4hkLxuxtlVN9AUKAzPD5XOlQYYswPp9gxhXxFgrRAJ8OGAh7pf7LWcq5giY
jMfY+o+dsyHI42hHaSm4eTfuAaj1aOVccFcLJlVfROw62VBnQJS4+oljIeXFRxZJsnXJVHfL1Nu4
qM2cSWw1krY2sgYPDOjtNwEL+ei2otUmgmFPW3UtuDYP6pQmcjG7cKQSYGKEc2c54marbircuolQ
yTjJcjt8kRm/ZFZPT2Yc2lhsE80N+ffjdrbVTY2pdp+owR8IjqUGxJxdeV6qQko1ey1LNEZrN/LF
pFE/WyOd8iXLK0JDM7EKAklNPo/+JOmT+stAsH5dymfxlfqIp11S5JqiSjKwUvzytcGobhbKk3k5
026ikr+hJTh5FzZymafx6NHRIjwCbk6OpxXw5XAGBn8jOMApOzl6CFlVQMz+oYbc5V7lUFAQRpDP
TySlKRN3nLcO5bJp26patQeHJe6GGP/Y/lOrJPkOJS/NR5+TBac1+KYnyPUq+Y6200oYzkLSkb9G
oirJv4u2aoUNOOiBx5aJIB03aOG313cnRAxeYz6y9TzRPgnKx5AJkShRt/SbKuNk7zYUIeQPy6RC
znbtB0lkXw8HrGnfqBfmcf3rK0SiWunkkPftzPYsxHr0Pf6Tuast9rTNJu2LRsbXPlYwMTubVCFm
a1Ap9wGbOMX/7Rcy5h8yvRN6W0jVSAiP5h+Af9zECXQmBqg9mEaR8Qj5OMgjveR0+5aJ/NFjcmfk
/J29cGw26y/4S2i4ls7wDC2omWnDU3bTM808hl4Js4RaIhel+vZMWH4tdEHIgIwex0gcgSZ2osgC
V2SbWYqvaE18u71Wf4/bDRAexOPZSqz+4lHk4VOq8Vgd7B4rFEKE+QmdHZQ65+zY8LtgZY8EK2lr
OrVn+AZ3XAR54W0EOzhuBvHKIFwEYLhSFjtGq5XGhxESrpkiZ35Q3rQo3OGGiXsC72UwyaHqOwdu
vWqmbO4Ycrh98ud4hxlKD7u9w9hmwY28teCCeDGsHoKDJ2OI0nFJtcmdwH+Al7NXf4JncuYsL9zv
z+dz6PlgJSrdg8YDE/ugWIyy1LeNZXlMq7Et/KRdbPqSY9kAulb2PpBDc6LBsBdmbgfx84Mlvv8D
dBmPcBOMaf32gaUdgar7CHHBGZPMm3Yx/a2JBpitVSMRoL3i/fFiVECtRZbt1/qPXdW9LdWRSP0Z
umQnkj07SFNYsnSQZzY8WQGO8RxJ/YO2iYGlhZRqcysBQDxLPZqNBms7yDR2180HKYiofp+mvs5T
tWbJrBl+Ap5SEngJa05kAKqvFeY/bikG5QXLp7+PHxoQ2Ls2u9fjp2WVXKwfFaAerI+yc+kMGI3P
mbNwQ+AvKnks6pmGo06+N1QckwcqNiNQ3kRfrKBgDvj4lSi3JnOz/Bpc/omt6nPINRrld0XtbBle
Ec8puNgUrx7UONVMccjlKyKmR+ZMiVmP9NMpd+JH8NVqf6vjnUxyos4Z7X6J393kdrPNLlGFgul5
J6RG9hUDLCucOhSuGfune72qDH7tH5q+FOMS3ea1VSBCgmKp+glXDJ8eUwdP3+jJLBU+PzeesDXj
xNbQDIKoz5wXdLdm92ujdERbY0VCmRKIvuAq0owq3eoi/TCwUm8PwB1x37XenZG9TvIbYJPWDj2h
tgNYArMkxDOt22eCShKXyJE2Uy3gvzOI6idJJ1+eVEV0hrqz+vV+HgBqola7uQOzQVEfJj7oHCBX
OpEd32zfR/d8PN0lMBvplozJT3BmsPU6837rrjeVoBjoZUyLS+55Y1j/VLlJqtM8shS1npEPAh01
WOH44cpDLLM6W8oruV0Qfj7Ur5Dt9B75CXRWVhp9/LNQ5KH8XtJK8eMyDM+GdT6b2N0ZFlp/8j65
unS32DUXMGk1nJVmjuZ19qw0gWHg2KW4LIdYNDIYky2ZRLriOhSoIZlCWnja+yhlzynhq6PYUtdj
X4JNTitEieDF9OmhDpkjDLx3w6RTClPGPQx9jelLHmGZK1aY2QGsUxzKQoFGVcv27cw717+NPc9M
4VoupiLylVU55kbtX4irdhOP10vhzB0xvRbnJDhgCB6cA57YU/7cTiNDFK1EIHLwJ4hLpyiUyWpz
okbCWmsiD6hawzVjtuniYP/+y7gLolA4JFo9wetjNYsKaPdLFEvjEnkPcioy8CHgm8Pem5wsX865
YOx/KPxHqIXnHBv8DhCfoqGu/6e/cFHCGaHFcd9YaIxh/DJ5+1eBEEUZywgWyCO7T1wx8Btw84r2
Px1eU67ebUc1vnXt3/8OHXvo1yucmI3cd0ODFm8zMinB+g98StoqPLce3kvx9K5v1U3ptQbJdQrV
q9XcwB1jflVcSi2x3/rcHZgdykSIizmlWRru9c2xf1kcS9gJF3c6T3MjYNAM0m6Mhp+fYIZsJOY+
wys5w0aEr4/gxcsVdBjEw5gk+2pDdcDn5RSdK0V0Lz2vF/6Cef3zkmI1OvHWbBAG7FL/HjBYSRur
ACTZzxv7fUPylhhHButVx4QqP6Gzcu+BB1xXcSWxm8XEejpogSQKn1Yh5TXtMLVFhMFboeX/D4HK
i7JXEQk8qul3HBCWEc9UKDhV8MeAvvdiFxPKMTxVW31wjVWsZAcCqqJUU8dzBBX5VejuGoJLxKiH
Pgsaup0Vf9Wpta4L/OdbVhuIYB9EbIv/cqDqcWiR9iAvH3iyIcS4RnM3V5NppPoi5IG/gSY2vP80
Qa5W8/lw8EC4tTk+xHhH+0UZR0Y7xSocTYRTbtQnQueC8kh99kT5Ef/N1yHYpuGYQ3rx0z3rBnUJ
6Ccp6YZjdZBbYYIrxWYHqx7nGNf9XJK1OIKZtCLkRs0uQI8q8iOSugXvaBJgjV0eBLMWpMDWNNsA
AKW/gsi3z+8zS59z1TbRsG7Pt5xQdoLGW2mzezdBr5nqJCf2yzbunrrXguo9i9KTZluae98AzruO
+P1S7GD8HikCcUxfSjbyutw6kv/HzHL1agEMBDFQM+JQZfKDjbJtWbVzSUD6bqkADVp5qKJ9+7EG
itr3jGLng7+ipjqmBE2RBMk+nKVp8+tLjxH55Fwfr0A6vygUndHSZhxv2YfQ0T8qV/rImQyOnPKZ
wqwPjCqGnowmbKQA+M0QbAqfYkU3p3AAXa7/2BtWbPftta/ffGz7Kh92+Mvfb2RAVWh2FwcVWQI8
0KAOF8+bFEmYj5a27OMGLVPM2zEH4mtw7pm9K5k0DAItDyKzqp43YjGp5wWhP7iqz3+eUrdwZJyl
ApcU+DY3bt6ktOfHJXFoRipqsKm8GsqbZyajAMyaLIVFuD2mtuAHuWX5t/aLBvtsPDiSVpk+d8Y0
YhywEpGA75VJBp8h015ZWCOFvT6fDjvH9YQh4hCsWZdNLQIeyoTUBzYNA7BNJNe2Yt+xVwiN9Irp
WoAasJlOBJdrqdpj8vP++87GwM7gEC62hcKrK4/IF/G0tYUZOtlPU4XmfFP3O+PH3svkTJgsb/Ai
Ceu7swBIYC1kNu7zErP7bwhkP0VH/SpO1qS/DpiJE1lspGy2cCUjIV+Yx5OgCacZONxlvn+G4Ko7
u4/zID3FRLau+grHIHyAfVNvWBEAZy4FadDSUC7ihupn/scv4eiIu6Ibu+ld9T0Box4ls3ntX2ji
KLdHWY0o8gUPGQ4fStQjavYTaQA5rvDG5Yt1069k+7p4dpNCfqDVIPkLlpuxmgO2ncIwhbrWye98
wkeTbpRTjnX+VAwmLGbZ8TwzF+d6OkeloGvjX3NbbMeQuXam77N/KUVkkyVQhVgi76REGfsYuCyq
NKUXxPkagkQcCAjc+MNOzljuIKm2YjA/vQf8Jx/5KrUru27V2DddLnWPs8gbF2LzBv6AWAuh0Hc+
6y7huPPUnBW0EZgr4g21MkPby683s/adY02ocgCDKRqasEqc4AgU11WKVQ1OG3YnWRhvh4RdlWv1
IdBNJu4AKFOUcKycJSxnjVb/AoS7dXex7QVU6LtiZb+zRUems+3YSG/4LPa4G61v60n4sOqRtY9r
JQ59rbxuOJ4NahXXW/r49OUdcP830EAEArMLJ7Cwz47xZMC2VOERv3pOOVCmmkyfXrOr/yrPNjG4
Vi7t7sQm3Ed5FZxIhd2dx4oG68KLMPNlB5SURA0sPuyY7hsGZaKteYahiFAe1galbyDKZ+DHOLM3
nSs2mBWWqYz1DPgkkGFWd6Ojfdew2MGuP8zo8w/qbZbM9DF4Dx4DA9dgVGzfJEpeBOMIOs+BRE0z
fb3veDDRT6Pt0hSffAjBG1abLWLOOg31ro5ZWzDHvoUPmJPDGb94kpxyvs1lLf1K7tlnxXcFr1Bu
k4lr2RdYWbcO/n94xk3/Upac8E13qZaptWHgH70UAna6EtikSK/Z+tb1JTYXUNAFqVaQgSvh2IQu
hhDqGThmzrLQb/6T1TZj+aVp9KuqYcN4GUcbtb3xLvoeLxm7LpeXXhIRi1bCvXqHmVUdi3RM57Qm
M1YoGRw0TxGP0i5h9jh5RdxLfHoCmgkVOQ9GMoU13Y9ZfimbKQ37TlEMeukBPjAxSa30RhYB3yvr
tf4vxSpXsLTfSWa7z8gWLQBNzTOXJ4UEimNQrHc9VMdzZrKrtuyYckI07UEdF7Oc+NlgeT4OOJVW
vDES7BuWyvKAncNeX54NX8fA2ClYvq9A6tmd9OX3/nB1rRRx33nfUYPSzaYhcMofA9qulLFEWUrS
WUsUP6slNmFfcM7ALHsF4AAhB3qyaz4NiM6IxjiRJHnXRx4O2bUIENtmKHMNYiTal+UZD07lA/Nv
jb3SxtXn79429+FLkbU67LKxoqxIUYX7A6oeoPhMFW4olLgkORx6U0RViLtFyiN8BY4cyR3c5DOE
WIfO8EeP/0m/l/hgl/6fnVdeQBHcCgqcPiHrApDaqnt1sIENs+Hr2cGZQ3XdUSheU2WvBOzE3gqC
4/PrqkDD67w9HbGEDGHT+hCtDY5LMnFZNnSq0q9MOhvKPt6kozU6y1PzVtaxjd58KTVzi2g14jt3
NIOgPKwRWc6KtGr9XfnxdJsEZ/+iPwVilE7r+i2zmcYOxJNHE6heDWf2Cohm05XRkZ8O9rLIIir4
npSebNj0lATfu9vxF0V7/xPC9jU5YauIDdqpH8nFO10S5iPUPTUje4o6wVBxIEB37+smam4F5/vd
8fUZjGWK/44rWokwAE5BzH3wOwdGjtEca2z8P/HJFzIoT19/3HMLmX3/MZdBSGZbEwOSbrUzNRSL
asPwQu6ru8iQeUJubTGF76GA0NgjTUiNvvYXNvP18ULe6gjjaYY5XGdvSGaSlkJVSRhUVqt9sNfv
8UaqHoVTKPw2vVn4Ygd8f002gU7TNXnv/hwg3nF2A6fBrvvru9uti4/ZIoQe3LpmGezsj3Ia4v3p
75pgOYMQ+fHcdAuAH7dRi9x+J9QzmBbHKALFIjoIYCJRBvaBz9p1juCPZij222HBmT/O0NUGUAg2
CZtDXJDDgrsM6kY3h2XiE+qVPu45GdT6bQ0n+GEEdQ68C01OUS0s4Y3JAFVULacSYJvaXAwGT6qc
Pwq4GzywIIGrr58tih9LUvX5b+j9eO0zB4ChmGxzTj8B/LZRenLVFDqNB5/DBwYg/gUHvo6+SmTd
uKj10Lcmab8jgBzsrzhc3ko6CwgsrevyOfrd/gO/R53jGYDEHHQWYlgGh/KmXSemSiXM+atKF2+o
52zcajLkMmg4Ms3jMQzO+26eohBzBtwRRIwqQgeYnXeA+pEBKCXvjXpTtvfz7U6wrHV4KBOGrpB0
BWrSGSQack/UgSw95WUjd5b0M0KvwKLHjKfq4qPQpvVLlRBxma3Z3OZSnhvrgM9dQFnuaWeF30vS
sAXwfJ9V0RNR9sUg4h8PnU0M7T6xgrxtYv25eyXUlLWWM/B4VhQq5Q2Ck00ENWMiZ4LjfSsioAkJ
nM9yBACGLSqyPa16AAIuqWQIPAGwf2y6dI7VR/cXb/6NNY9ih7wD0KqDXHXg1nAGz4r8GSIi0hP4
K20Nxq7Cy7Uk0wqyxq0PEsMmnGl3wU3vsD/1PPvIbv+kT3FryQY5UiO6CJ0GH9fn8g1RkoRk8x++
gp8ROOORhjUG3aZ/zCEk0C4patvjxVbqDA1mDCtjRVxzEErMzV+xlldeH+TJvP1QlSyP+9XCPtTL
zypq2lK/bUazINu3BPmsN5DHwk989KNceGA4bt7FDbncUUF3iX9ALFExJvHgJGP2AeO3XUFje+Mm
iehBsVN8gm/XXP2FY6I5rzdEggDAXho67CCmVUoV2qtgX1iI3DIO+iBGPkyW463wCujnc8oC4zE7
gb3G+hU2FjkQoSXcz1hVHkbee6QZnqYpT5/oKVQPXRGJ5lSd3NN7VbDWxj0tvnyrFhyV63U/ujJ1
+yewk5iOkbKy2yQJDBLfgcnujTsb13OBtdxcGJ/ucIhONtojW73AdmhQ5Q0aebbhOmRIyLuW0Irj
Dad9Mhly8W0ioRMYyw/nDXcSLO01Ob4M4iQT1bQ7v7PFZC0X2BVbOZVl5zobrxReOV8Dq4nBRL1F
8os64yQJSXyvJZ6mv0ZXGeyoDkV4C9YW3nSnkhJNFQjv0H8jPxdmiidLyWzDEaYYbzOQ8XzgIrQj
tLitfBgzY7xe4jaCWw32AoUkYQwiBQbJMXvYigg/VGAwoCseZse+OGGWfdDC4Sv+RXCXqeNBpdOK
Jt9+H6vZizyWjj5Oks1S7mL+6/1m3R2ppA+7vi0iQ7Cz0Ndh1FQzmAIr8nCzgDjka7YqMfEwZ5Es
n/3wgnz0LKDHLRMyOGyGLH0d2k/HOY94G/fr4bFAt0hjsOZ+HZ0+YYAdC6UIjZUvCBNS7beoLiwZ
Qs0AqBWlvJ3a6LfWBcjoxCcuww+cOO8tXKniwqe7IAbxSTn4Xr6/DlZV/WuRrunMqaYbfOI2nqiw
JOVS116ivEsSiaC9jRW55aRPF3tOa8aXDc+XKLagf69nOAvkFWzWHNzTxy4qYxQiNSmXRZGAkXoE
aeqNBdJskaFvC62ooLiuDT+e6mnAe29xgd+isgkB9mhwdWYwPaSI02PblygTeq1LBMgAh8G1B9TS
MTRYwFpnfSji+BbMG5bSZ5EId5HPT2QYIthTqjYHICutGCp2zGR+wpk8Tsbkv7e4AIkYbgaWshGd
zix7LuenjNgsuCXt2tU0SBCOHcyDl739y5PNX42xLJkAskrMFOa2KFviYHOQq+fMiFF3l6yOtHr8
ZCnb2T+7dszhVnT33mkAWzrRBBqg0kwxv5Zs2UsEuR8cN1qjRo7Wf2kaW4s6cGQlLK39J5oRv2sa
7MGxMpeEH9rp8e8ChZSOEhcgucR2FPR4EFo+lq4Px6yfMWcjtEh6Sn68RCbDadX0iYksCTaOvk/E
ZwfuNZx4+yxgpeSmdvgTzz/Pf6mO2SahaTTLXvK0rPpFWIElUOyYUJ27+vmykzZ0bjEYqTT/WS6A
BvNvK8z0LoNPkW25zD/BrIu84vUox9+wbNE2VtN67dzc8hVFHBmZFjeXaNftSuCp6t/+o7cHBkWD
e5QkTSDxKAq+V9BPw8WnxlYGTE6xnYJNRGEBkul8zBAgvCftKUwKoKRi/lyCBSTMRYU/rzUXGt+A
YGmSdvglk8X5v8/VgnbHU/yj2cr2XqIbMqTnJKJVBeLDF2f7tk4wU+A+hrg6tAWmpIDGX7kqil/g
FmpeX0lroT+6rBBoKk092xXsRsZj7G99VRCJQAl3gFC5bBBhzIsNrySTFL0NtSsy4laoUm6Zb4KV
BDTUW1qryXQvuK3rFO5Jy5LnX2j8yKAkhL7KKRcvi17byX16lbAyMbkcn5E6xUzTftBn5QLbqyK4
QiLI+5UwUXtDoXkjT53kTLKXQaa/QR3TtbPRybgrIVMAjuyXARivTDcKiSc9tX+5F/CVdULhVkYf
3u2LYtHEqQZSa4OYHm5RQoLEMllleR/zhupg21Z+ofplMgoesRKcHvn0nI5JBJdU9xZ0Ihw1PPpb
Z1EaTDk+bPGUhWO4jOlUHnDRsdpjiR9fyHUMjRM2zZ5DD+mpSrSpw46GI9BOV7tnGBkKSscpjbUt
eHPwQbeUhn7fJey2VKiXAy0CSHOE91pRzx64ec4f5+Lb3jYE7ugfw3jB974sYLthNQqzBm2zYUiq
kX6UhuO8LZfkjr9G8ZGR9kGqXxrSNOAV4MLzvp2YKsqGKblMboqyqMWMFWNTOH6jrG7ScYx8y6Mp
oqoYO4vqH3jEVHU9+ZhA4i1OEYRvssKRI5IRp+xB858bWSO/azhax852XZ4TmXaUyJvJNwzgn61N
mnRnMC64YcdUQC+/UIheKvBwlhJop1R2q4qgndrZilOFrEX2bNB0FYocb4Uj758B+ZbesVNtgPGp
2GsWsP5BuetkZIeQOxYdToYEFxA0dtCSKhWS9bMfHM6EYImhuigbRwbvnfYLoyvS9+ZgmFKe0CG0
d5GlgbV9Ndbs2NX3rzIAjLzINFqgQbqTooX8KeQ+lXsxFrMXyyt9QIyTZcQ66kXJoKEJJgq5bNeF
y9zvW0RX0AjEJy1DDqS3v8MZ8xPBBvTjSbOBYf8crS+w1RO5TrGNKT44Aln4R2ThcaXwJ7sYzVGj
viDZa4MNfswgzYUaFppqP+l5IliQTkbuUqfzORWBnH7KS3mgAN7vJRaywl0wAMD+0KCMX/xppuwR
r+JUZSuBr7MLQ5dI+6BmxwL30euvQe1tAvgvz2DghBV8JkOdX7OzXc5IaGeUf4IwKWn92fXWnwnJ
ilTvxJwWQm6aA+x0ISGfzo2rmFGR0/WDTzNtYazvt25BsDpMyEjnlWaGHa3egF5JkjHh3EBjsJdZ
AlxpA0hQn1dt7FXWZStCt8f4UV068AYABFaRQ/DHShakriCg1LnQ8L3Z8+GaS3AyfVfO7Ut+zHnQ
bTS8/FdUJPxCIhvoXDcBp90wmsVolTeGrk8KGtYTbe37m+IAJt8cyq4k/SkxWfWeBVqhj0diu3cy
5ydRqrgLWACknlpaYkr5gzMBpFvGfNY4GM226hb1NdHKDVvL1/VTsQ4NCXhuHZInt/k5J2Si2fdK
NoPDk7pC8gBxvgypNLxeSsieCkptx78EZFYQd/WtDILI/radUGmFyHFxGAp8M7ileMO3BwrHqskd
XVbhbrQTgCIkWxyUbWx/OWTTxsZsFSHKRANsUrMIf+gXVYeJVmuHtkNJ3jUaum/YCngbDU2IcRrL
0BGreybfGmCObV/Y2NjXapjL1oe1YmZeR/H0GmK831Ws3DggIgu4gA7MGFakDR76CJl+mJcCJyCI
RHDFji43COEMbGVxSx486CofRmVdX8ZiAvuF+Qzt0ohsH7uxVaHwFdViC1UHjsmE4aK919SVxuAn
ganvqy5f+Tq1oyA8MTpeopKiocZ5CBHE4BcVSy6IrF0WS7fEUEOzrSvT4cylvy+1YmXxsN5ALqQh
cgaV0bVW532H6+l/Wl0ac1+Egg7I6C5oU8ncvFmAa9/NfTu7sFYwrNiZsOb86UxEUnan484wAo+u
IzjflYIqygvQpWqx0Q1cMfBfIIiO4YOgIrtCp4jDfQTNUXegEdCJI4Q1qHVmECTuK9W+PQx2bE/o
5EB3Ute3yQkNiZg4ZqwhPUQiM4PFLj1i4Y5XBsgJphgb7w9Vz3DwVnYuvUd7KEVNA8S78/xhz1ey
CcQdjNCjwAdtW3O0kPxinx8NiNW7dkIBy3kJaidTzA3+ezqwnYmBBFAotYrZLCDYeYAUEl97o1GL
rp3LXcVMUrMDl16cWG+vaEC0m9Hn86PXglN9xA+u+lMwyIzfZeVsuDfYvWNe274eQ9AHy+ILFFzJ
IlsCO+L+Sq15/PPSgIHxmDxYGgoqg54V9V1gNB8Xh1S8e63bmDVnQTuvUxoDci2/bdlE8j6w2lub
Q7CnOFVzXg2d/zz7y6iKZq+2DXjOri7HuVQ1gHajwTvTpb4EpZcl552B0St6LyUaPli0mOq9H5U9
0QJ+UKY7IImtJM0oDZ/yQZUdHGgGCb4B1X7DpHqQVJbYPcyX4Hdzk8Udz6Zw3iQIv6c3a8bQ4BVH
kxTGaES8SidmIujwefh9G4o9RLOUBNyKmNdc4fYCx8GKS0LGvwuYRANsPvFM4VNJ/8BPzuStDG/0
2Et4Idkd+8VAP02RRGBBBMy25fJwzM+P+nJRa23Ep9Fz1K5uvfm/bG+YKID9rIjdZZ5Tn6Qi1cJK
6kkM6Rxu8x0FkiB7Ovmi8SwtpyCetVOG5hY7zYPgkv4imnJPfG0e7BRmXVBYNBaY6opLL5W4zAEZ
N182xqcLvzSAdU5giFfyeS1VEwtzmETxfqjHExWrBWqj64lznmiPWSXYsv2wVGpfKCTgTOobUKF6
BaGsdvnLXsmlMCj6tB3/O1MAQXzPvtmQcpWPVmS6Eqxk3O9QJKcaDud4mfeZzzfsXZ2TB9xYB0Ls
g/SolQxMwK5OFd5sPdJ9etQaYJm8pxDJJ6Pzr8nyN0iIiqf3FI0i9EUyiW3f5wI0diwu8IHF3RMu
b9YVglUvZFtlppiUSuLjX++OIcxw8JJncZDllr7kKfx4gfLtsGtqtX01ShP8hvFWxcb47vO/h7zl
nwXQ2zPkItPo8K4TScNBa8xpYINULs4RY1ujKuBkSb2eBRFhZ/R9B0cJAVYg61bemym3Kcokjxm4
ieR6HePdT7B71Yl1Ipu/aIIdc+YHfvMb/YEDAjct0UtwzS2AWSY4I2swHVRjLMexz4hDDvciARfg
fBYXy7j2SnvnuWN0ZZAe37XQhXh6iOE+/gOBV6JnAPGBj63R7bH9+kJx21yQIEVsaQ15/+RqBVNK
mqU79jJM1cQF+ibRnsv0wuqJh4eSCbFfyIntT/r0ttu6dypslvuxpEWV5eWs/0+h0zhA+1gJSB/k
a3O95+K+/KqY6ifzPVS4MnkrFhR1eYbve/6ERIQa+NXNjza3TldqusNufPWVacItigKbOEIsbpsM
65wWfJWP6n4TW2XkjtD7se+eU7SRmoG1S6660FaZw2fNH79C4H8WWo+SFwEzIGZdSj9vG9HEH7Ic
GstRcVtzxsaP3fM1dlS5O9jZp2fMbaUl6Pb4aEApCXXkKTFoHW6PcvtNMSWnXTpFgj2SMdf0hgNu
cxhiI+XKsKMK21fE6Z1FSCDYGwne182aoS5yE3j3BZs5rmMVhRH4+bKexRFpAffliiHnZP9ilEIS
vXgOcQxO7Pgk3VNeGkotLPHk2mKH/u6UKe616CWjXvARoPjg3A6yjM/i67uePFszFXsXzaB+4S5j
BBgIQ4Ikg6HFHH5y/NBVwzKjNwOGfSoMwcgrzIiwAkbmw+jV/HbVNBAMaqcQVOtKfqqjHrUtu+Zr
aoj3ZPz3wxvLwdhWrjyq21hgrYmn1RGT5Y6l82MW5vGEMTRakLTpd97sEy4n8r5aenoFl3w6DJXX
muXprSKdCydRffN8/BEI8369HiyFEWfu207iSN0Adl4NCHCLMVihG+dFZSZJupifla4eJXTOF0lY
NhcZVjyxHjv6jJcQ+bdhM3i4Bb1NM4Crppq+WUlgA6uCeXWSHFFZzn9WR3vgf1gTo8th6WT+Qw1Z
wpXEp7/Sf/1XgdiKr3DiRYm/coVQOx62xKLrYchzHyil3FXPzIG+eBYUdlvx6XbitMnAWaBLdB0d
l5mpQoyJBK/+35augVlldLuHKZjp++HrNWgBXztlOIXMykbi6F3BC6+7Q1+KnUnFYXKhrVF29lg8
V2lYj78XaEUK5lqdlCc1rNeFHfvFAJkWzidjDqcl/Qp2Htj8q+NjHvn7Cr9cFjkNxclmiorAH5yE
zSl1CDLjVjdxL3iC5IZt21FsBIe6Odhdy6he+ablWYS4zZTY20UsbkPfTt3tyN+C20mNnGRVvvwr
eO0hluxU9d8OM+Q9GxFhSCOxJmoTvdft0Z7CxRR0hnEHHzvG62D63JyRJjC8LaaOrUpCQYX21Td+
AeZxvNVTmpUDrTlUtY43lXfJszIDoYfBaaNkS284LERs94V3IQwqDGRgJXByNdd3k3nHtCLc/VEb
GgLYUG4z5lYmc6x0xiSdnnZzy+8GotF0c+fxQxnLDSF3aPLgWWNajnmCYmoyncdZsvwEhrX7NWnZ
4ylh+jMDOap8iMORDjDYgbMTESEtm/SyFI2PRb3jHczED86f1KQOCSu6dT1Cpeeo2HYISwA26RkS
CuqutRVtGribzP636RGG4fXW4A/Ao0leVYRIJ4BFbA0NjFjjzjlOa+qEOK8R5wmn6lwI+wH80bD1
O2tEI9aw6N80iEudI8MLUvof3Zte5m+pYKuRf0yyCJ7N7z2qRJ63Jt5JZIPPM9NLFvEYbVk9Ryg2
BjsYkokY5qxYKMCKfCxlHOzCTPsGB3pprIPpCUH2yw7KlkEwcBKkgnIOnISbDyx5zYQy1bZWS91w
lQV9SxkRbtWeAXlmna/nv1z6KJpJUPmX3QFuy2PEK0rZnOFf+/N7UfBpyD+87LAUDxGNfnVoimNs
e9n9/wnURQEy39q5GNihfZ6zdvVcD6gHiYFk1BtZ08e6iF/YbvRviRFjExT8O2kMvApKqE9nZPKd
PcyyKGNECPFCMdVgx+rg7AcXc96vzi+IQ54LkbSBloGfEJYjqzW5VqnqBZ+aOSPwiw/qFXjLx5HO
c9tr0MjydlHlpxJDu+HXUaFusjEerM3cSSNfMU/+QEjk0C040MUyeKDha8RxDdp7l+n9p4w1YMKn
lLv16dblTQ0jjjIp01BQOJ2izbztJwjfqN0L2zMnMu9dTtZI2Pwt/6MDoG8UY2S7ic6a3IxomSnx
8J1lzFgQ2ZQfVyrt02WRywOzCQkknx5JsOveQSl3+ooZJmmQEVA3nq85HWka6A5+cw6IIfSa8jMT
LOFxThfvVkAVNbutJfKURzENlScLF9gBMzT4YcWfEbBXY8IA8F2qyd+IiIJwnHou72L3dP+QJECT
Y+84L6KCByLhLUkjM6HsnzJWNyIUgM9+AN4CYMm3WgYy8KqEp6QqQORg8ErsTAjWahKmGOdwkvzK
0TH/5yQ0fBJG9qtb0SSquCoSTSpNtlsSH9WlAroJ/bq93e2hTCIMF/+Y64wodCo4Q5RJBrIiRY2k
KN0Re8n58ANKnCJj4NfXPztPvfTxWWtrOQ/z2y1JPXNBsS/P1zIwVAfQiks9ZSFWhHkBitOHldFE
6goyHQOFrHTMO2ic+ei7GvAoCXWAHlNOs8zdVSWe32b0RB2OYZhknBnCfogixvVNhs3zfmALO64Z
8xC+z8TSPKUAF73ZXdpn0vVv9yDJbzIaggylbp5txeIMqe1uQxRs+d2XNJo/+U4MWJZUKuYMbk6C
VNhKINnWuZ+a21sLCjBw+1SR93BrI/WZkzLM6UGTnJFWEbMFvy3JefamwIP2C3aICVQ7cJN3BwN1
MLlHxRuH0hxfabUjUU8W0qrYDaobeeTwZA4cBp6R2GpYPQ7aPnTVm+nKOXvqcXNKsgg3Hhv+7aeO
lMLPYWat5c9vn/ldlb9k5cPtgUvYMPZbEPPUCwBzofTziCl54Ch0DIeOe/0ePr4IrDcrge6todpo
HBgkTMSoMK5HHEkHuYmUscCg3lY3Mgk7aZki9oX2Q382CDvc7P5ephWoRj7EZWpPCdlfnMRWA+Pv
wf32rfNJWqMv2UDeqajDgmHdf54pLmbXDT+Q9sVHhZLuueee7IE5hizoFB7saBw8NKDtSnhmNGrS
aNq0+u9y2vo1WUDloldDuh/VOcmruNaNy57eWm7RzY3w06fdOqDzJ+IJN23RD0QpkPsHDF4us285
00g98Gll67qLyoIpmvQ61GDP5EbIjGViw79Y3ffkZ0nqR3TSBV1mYEaFqhy2PA3BnM6WSzVVI6tC
yQYKf8RkD4nlnK1unP0lz7yeM956HYSte2DW0hITvDVqhPnfr6bhkYkQ96lbIgUjI15jrZFk+VUO
Cu01E9+nA4+DhNcRzKVqyn7ZyBluuyVPrxagPBJIl3y/u8tTrsxR4igFTRaCRCPkMWDk7eUfCzhy
Sc07/aiIjXpx0dtB0hsRxnQxflOQYjO9L0B0CzAQWsfAfPTr9Ne3V/xBtJIm0FhEY3jgVGYbRuL3
n9AF4MrRpHH0bnAH3bkso9S2fNUeLhhz737wEtUWcih7xZ+tMiXvZir4AcXTSUJO+Zgr3KPCW2ws
gmj17Pf7iHxTfgVE+5VNbUCsJhKFifhGoNajnTRLyaCZecuBLSQFzmvPOqM3l+Kva4EWRKtFaFwG
JpjPRBG5FDJ4kzWeu7jmiRUPPp+xpAhu7jFKhJ0CseNb7Yy/WCkPtvS20LhyC2bEmQNXzqQLX69i
M83NKxpaIqRZLk6T1IHjPgLf2YQD5mTiuFdGOBO7+HsIs+Fyxvh9B8XM9Ye8NQcSUE3JX3kQ2WZP
9L24qKWq2ppbLgux7PXGxJohFoPId2HRRzSwYeizT14lqin6KBlRROUk7xtifpE/knVPtAKu2lw2
QPoYznnoB0aAC6iKUjFpYx0jQlcgwHlP/XpkYq8DU4BgxtSD1d3nudHKPpMQ0uC149oOfiRSRStk
Gi1En3WDbyCLJcLXULz6cq19XZYYqC3uRp74QV52QOquzyave1qJSQ0sdQ4LfRCbk3lsmzQCbwX6
qtj6YLAxrNNnLohG8s9/e2h0u0EgUz+Sz0zkkcIgBXmpue721XIvq2DDqrsJhzoBeLU+ivmqjiiZ
akmzjRixXo49HTOa8SEyO643HV5Ft2D70rXkzoYob8R2gFIYM3dApbbDg3W6yfWp7gGXKKbbtWK7
Ot5dNG93g3FHr33cMcEpYzGNK1qyZYrdaMFh/08kzzlkqRWY7tnc/szgVjqtPH1dXKudlqrRvGtw
FgHIblUWaKyoZG0DBossJ37xnvcWW+XUG8vw62YEbC3vmfEyn9K7PoS0DwZyIbUsGRCrlO1fth8M
ndsCiT2K1I6bPi0iK2rg4YqBiz1B8tzC75RXir4Hdfpv84eQ4guC8LfwZFLhQfHuPqrHjZmzkFUD
fKhEfTYJknjO4z/Ohka0nRtdWfHtt7Nob3EpGbaEF535TvkVqqFNtlNp7HzNW3mScexYZnCZmovy
6ZtEsih5sdjpsevSRQD8BYv4cZdlK4FDXuFG+tsDWlO5nceaAuGxTBc9hAAM2HhOqbdjEWP3GMFE
v98V9As/auGYPOgRNpv4YBtrq6ggGOjLEy6hmIRTtD4EykUeaq6WX31HRwiGVm64p4Rw9fu8xeHZ
26ZiGhBprWj73UDfuhd4CfGccWP12usKtwwHl+s4+oefHuZ3L9UvgZHAuN8GfPC+klgx6yWyJXTH
kPoVHnSkxVo/STlDPVDadTkw+RK2iejxfntbBAj8jqv8r1TZL8HMtR/+wEwfrnjS+m0SfchnFcEK
rBfK2T2yQe+yYWaIPFquRJwxK3H0870728hHFkdbQ7eSL7V/6TpDqYdMk37aSwkor19VghbCqxSE
X5+XQhn2sJcLJp7iELbAxWGn0CU18Vi/0fgdcFgmaqBUQrisonX6PuA7YIbyV1XADeh4J8U7VHN4
cbn5mfVax8ZjV05LYmKCLqzMRoalPbqWaXv2N7yvMGVWq2kaRL9br9OHzZmGihu/GwvSBlM7jOk2
r+G5ZHnvrTq/v97SWZmlLqvx8ZSZAt32bay0fkdbDeemGlb3sPsHAAdtLpciE91yKhMypoeg/Nef
VfFfgea0ia0SwRfP/Y5l4Q7NRuc7ejm1PCRCrQP6A1mWLcmVPzplk7PSY4RgtlMYNiD1Exv3lUeU
8zh1Tg5w8nSmHRIlwShoyo+Bbw/2XSt28fPlt/nyTLh97C1nj+2jmEu6kssjgGRhUyZsKoWlppEy
Gra9hTOZtpVYH/KnY0tVGj5cO3M0Vyea8Tqx7PRG2OecthBPqVYmerhNJbs/56UnqeQ6c0NJFe/D
lamE0t6ypP5PnE15NeA0CTp/C15GjXlTqpddv/6Hm8kBsHkrGkhDskSHmIgxxdfLEx32Tiy9VRiP
hhq115Igtdh9v6ytbz0zOAeS+y3rD+7JqBqfZDslbx83RJiTlJxaH9nZlmnj1A5RdhM9hOrGzKE7
pL+OKo0wPUw12+UizX3ZxeOaRlFWQbV11Hv4kTg55G6RS0pzWgfAAZC8EQcY2OXD4RRo98JihAIX
l2TM4FlPmcb8narEmpmkJ2P4QktlPDHjkSBknanicFbHFKgEvF3uleDf7mZ/7gy71r2nohwT45Qj
3waS3yoZMfkmlCYviSarTnmv6N3LCI20SjHV3+48DQHejLidoCtUu7dJGZKQMpw8ZeUMkXEFMwmA
aS22f5hOE9ZnIC9F4S5P7Q93yMPoMatdfHpGsQ4WJ14P8dXOx8R8L/NMPCKr+pfLuaSJZrRFSCBG
t2MCJmZNrcTGMqX8wvAWMVqd9CcNg1toKC5Snp3G8P+wS2Kbt0HTJSMpIC7swm3wkML4VyHbwUeX
wDqBDNTBA4YxdUBzD9GYIFTR1cH4DRg3/QLSax1q64tiE03NgwGrjXsdWIMeRiyiQSXj46u1UDN/
Ed9tdURGq64hTS4YwmIfoZViWAK1F7Oe23KROoHBv0ExvUEhH32YWfEIDos7CKvNYu3phxq+BL7F
mVeiqVrzSvaImIuCByMpThr10nqJiIRkucnMs96pFi71/BsIZU1fs/OVYh+gUJpxEAjYM5FywWmR
LmaH3RjD1cHjzYlHEb8j1KSX+cGU8wMXDyYhiqN8WmeuubwHhiihZ/Shr0ectuoe9yAP/BPi7kJJ
YiTHbqjQq30r4FoZXze7Yi6oSu+WnTWghyyW0uDqoKYBlceaHNoHG/QbbePga7Aspc1+YpvrBD0r
w+MWJxtpZlhc4gKQ0ut0qG2R2w0UA7Y0l7OdnagiTGjMtWkokDmGe3b6r97q+ZPWHLfHMok6Ki+s
N38A0iEy0JbEr1xbmKBhSFWwLE0Pu2MLF8N8Rlu45/imAXt6YpfkRLyQJp2DvH1Y1lkT0SCbRmhD
vFNCwd9YdyQRN5PQ6xPLsGzVslXJa0YDsQusMvvjcd10jLVZ7JaHvktOBCBAGX1Vn1jAmF/GFT5c
dHDOQZFczVsHJR33mQavHm+3QC4Pr3qghvPLKk1Ko0C1AlFA+vRvxZzNa8YDbv6O0fnz45DBdKDi
IdbK7UfAshfopNl+CxsIwyLcU0NZnxWDELAVzdfsFxE7jepqOM2P3+ozJI1IXuBfqy8AVI2TUWZv
/tjKd3u4xuCa+a2OVhW6j70W8Zt28g8TPG7UIsvRAcJ33nwXhHZpKgk5lvX4vetoeX0QdPol7WZy
GL1E7vgG5wVC7TXFfJQNTQcaubIutca3YfSI75iu+6tdXg4lYNRrfV9rhPsmuz+lfXKdtlX4k1+p
riND7747XxTaXMzV0hBkts6aySVIHK33XJSEPteTF234U9XSuhcubSwLCPS2joGb/Swf9FKapPK3
V5ADjluF6eO5uPrOljIEqgdDSRokcSNRETfK2TFxbcZ4JA26cKo2X5UGwZSXgici7Q2g/1BWb5QY
tFv+L2Mv3yulRdzvKe6M8Azd5ODErck8pNVOZkNln+vEULYEB0GcHiwAe6DgrslAA9vxocTs0vDW
BzSNd0Wn3zu5rVXPtMKH9gOkkmGIwpNf4pIIFJy9ZN776s+FPGNRHmDvGn2Nc2feDr9pQtJkSsDS
MkmFaZkKjEoEjrzaDStD7R/nozvzboUzknaKyRccksGNpv8hr3OgoPW7blVIdB4P0HCZ8UJwVlRF
jO0a5QHPJMD2yIoaxnu3JQ/QoIn1elNlpBs4UGsOvDTbTCDI6lcunKb8/XId5l2pfTvBnSM8b5ru
kWfu3v/VsRKuDw51wsWBWtxI4jQ/vodZb7LUS0Mv8ynqfEdlPogJfLvFiRrxwsSPBc0c5eEOtOLN
t0kvNS5HwqGtD3pqg8pe6yi5eNuXv5JQBJHw5t83ysHjvJArcjx8qOSygSSe2yExszW20GQWGXG8
kFSX0S88jvxEYeZf5IFHjNAcbCLqj/ICJw+Hc2+A51MUxlxWut9LziixVMzCvGDyN6HoOR+GRKts
zmGk2sv9WhhuEX6Ib1swfDIWkujoPcSqwIxwK6pabFAJLOJKv1M2tgTfiBiqSiT1jllfCQJIjCGQ
6vD/57vGg4Zo4Ea5fjcQwl1Ukn9bMeUxLJtoj+ub17OUOmrASPxyci13UkFoFAXBbUcfe63TxBtE
80f9k3Yt5TuLF2Vfhjm1r0j+FbBlUpyDqpNwI3vZYULCeel1Oec8Wmjm4LKIoFfW+4YrcR2Wgc1/
Nt1POwv7IlzweekDvR7CQqrfoKIb7gaz7bJrXMj0K4W3PG1ltYHQua7sF/XIXli6KjGNnbxLZ17g
jv69HRDQu4AejZ2A8/5z0R1SAFvlZ/dauCCS2TW0dpvKDYQQIHe97mD6V2Cizh83oezqa14AE7G0
ia9cjp35RbvaVnCEcn98d7RVfqh8Mcrc6ZmQ2u5SusqkZnNnJMPwhDYP79iFXqIOfWF78iKG2Hzi
eL1X2oXgYlWT+pJrVxjmBr4JLKJ8xhGULDvS+LJbwOdTINP55DL8d56+o02V4qb2a9atEkrUpqe4
mpGhBG7B3Hk8CrojXQyAQToHGI7INYxdfJ9mkd/ScvZ76HWwGzpd5pM6X6vIDy4IAUidEewHpGOh
wZHQ22m6rEIBfbRreQ4+vYeBn1wpNM4wMswn3acr3Xlgm2K/wflo0Qf72aiMGYYHMMB/NQ6/Fl0s
xlpKq5H1UeeMJSfZ6duTSfYMsaIjB+lkg49Resv0HziT/nJEp32cK8QI0lWGojbi5VJDZ2nfe3Ny
hNfvaMbnQMUgP+sJFPcliyHzmBkDA58ycLsyBghO/YBXGzffsWhEDCiNuIlEpJvT0VtHjZHQF2c9
Kqn77lTPqilDuGzDdibsqPacn2QsB5ra/hMLLah4KlqBhR7F5jLRGv5xHZI2WE6lTksJVbLLfTwc
k0kjISxA9+nvB/qhjxE/xZ8VggTJe2JvpsHli/ci+tTKGy5Dc3xW0/UCTmzFI0KjRwf5M/oMnVgK
L49VlM4PwzboUivivxydtobrRInqqB1tC3HYwwpF1T3PrqEd1FkCNbP3zzauV4spU9UFIwKCuEm5
2RWbMYKVVMJD0JraLP6xMlMLAjC6GDPl9l6th3/qkkrTSosgxgXMH5AXJ5kU0Lbp/hNinpveDUU8
V5QPP/QzQo9G84na3dUyQlNs9+pOhLDUo86n9DgriPrK0wu8r/WtaXCXNMkaQYm5dYPL66sgJ6Ao
0HTMDEqEqSWQ4oArhUoRSp7imz9LdRdtR597vpL3jcpRcFuih1hAo+Dd/0Uh7ySQSCodJYDO8NVF
w3zpgi3cfHrY5jZdjnSH0IjeUngj5EAjuDJM1wFrA2EZb1kXlyPyAlb017o53HCqx/txN49E92+E
t2Bnz8zbC2KEp9lG8pl1rT+m39ldcscyzZOU36zwn8ljzYGcyQqzrK67vjP7geWbLfWwByCV1yI9
832r9Oio8m9XHrG3OVWuNlViFQ6eGG7AvQd+XJVh28C/pPX9FAUAmOJYmM1IpRFk9iifzHVGcTKD
bz0tS0xvOgRoFfQ91ktaN+8TWtWYInTaFsIlQGyNJMpvSO0RoeXLfV8UGkl56v6JL49BhVdK0NKS
VP6vunI+sTRxm9irrFAoFDOPtjYu7o640LcjSYMA1Mne3jkMOLex+f2b/LinsgjsL89oXIajvtLG
coNfBxzu7xWunyc5DAfcjXUGWD1hLwtMJDk+jr2bDwx8nF2OVplsV/zx6cg6R7xl4mfDkGq1XYia
OVwyqCK6YEL/vo4ghEgiLvYcSVuIxOiWj/plO0voHsRX81Vbjsmr9q2S9ks/KUo5F8Wo1jnsVaM+
Kc2onQJxTmwzWTdEChrRu8JlVfS7b28qy3JMcw+LTd9Jr1gHeU/hLGJCbsqdoO7YDXpniOKQ4+tn
6TxvIKJnM9yF/B/vn4MNB+zUx0CEXg3ZuWiDcJ6p2Uo0Trv3WG3XCKqcpLFsFpTNNfBEcueVmLKu
6jUIrZDz3O1zfPGmdnE/oYW6e0uga46n2FeWL2/QD/nxkDCIfND3aQCD1aO/9bnmByH7ClpZP/0t
Gxd2pqzbXLUMQqiGVrrXnDU4LcKCcQ5Kz+AbXt742jiGXpMJWY0El9dnJMZKZ3umeb4Zm1Amjvb9
6K196YgkIjccqdf1gbA5UdeEshBjEGzs/ISNKnDdVKJzaP9UVHx4EU/vRyur5SrznFbDuC6QE7Qv
TS70wOsXbeSXphS6+olM0moumG3MjtpJTJjVk7MlDpUCcRu5x3Qrqvt2dkcdKsMcgUP546gkDxgG
vQ6weiG36WqYw1yoogfu382YtgQG9tUR477QPLPzWdlnmuDHXymiR5DhRxMTeiL69z5Zyk33tIzR
6LQ/m9/J3sraCkRpDgUQwoYucq+06hZ3xYk4DTl09huqrdN5It8lY6qB4w29ovqno+o7BRA67KZ5
K5n/B9tl1L4vp8uvpN0K5o92YV3xqGS363Dz2/DSJOCoBF8Ni7Y6OoJmJ4vnmovKn6c1PU8i5qEx
zT7f4agN4T9N+4BKQVLcQbHJt8nBk7jL/RDsf2ootWmcQoPL0FMHfZIu500/nbJXuhA9p4rckeSv
xQMc8aKBpeFRMyt+5ZKA6Jfn3KxUIH3R7iWi/8xYjSUTeVGWJ2p0qGcgDJE18chSP6bbsHGyMmWm
qHYl4H8ssbsHlS4aIorZjpPRm5sTfgqMUk3AOFl8pz7tZ+7MMZlGW+qFoaNJdd0/VML7v5wX/l3I
3G07xK1gxSmhKCbCUAq/hLLnu+34j2LjrX/vDMeg1XQO1mbY2jwXzYkdFKeC+3jrvXHl/hhSzgkE
Nkp0CFOfnk/6OO7HvSCORh52b/xHDjIqeYN1oGfOsdygBbqpyzRfJZ0ll/RTC0M3isyTyZZ6MJlS
nD11Fn0H8VEF+u/LdAcZnmEnidSPia86Zl63rFc29K7kjSAcDpZLJzbOiJ9V9vfgw7DvbdIlqCb9
cOGtdvC6ENFV/sd9t/KsR7h5AtyJsaCPSS08AyfFf7UAzzvYC7mtmVGrz9o2Ra9/cx/Ulur2fxyW
1TWBN04ZAK/t+MujVaSbByqcuKdXn9QC9flpSI6bkiyEbP93MWtaw+STMcu8Qh9Miq+1loEv18Ae
WVmkWMnvmYj9ROVuJTMRKXFej+6AopgxtBq5XJssn4VrGeQZQF9KK8ESX3bSaUkecx6s57IDmqNd
RJPz+13kTZW37q1g5VKtY7HU5yZf9Bgn3JR8K8QnoeCUaioYU6u7KTCvtH51rgJy2xL4zvoWUiP6
dfX+/Vd0lHvernD/XvN/ULfYGynD1FET+WM0Z/sRQx5g4M73T4HGTZQcOu7CiY5Dno1kjTW606S9
5dZ0P6sjP/CMWCOctLAb2/aO7n/V/lgp0RDD/XJdhRWhJaYAFme1bsDInyDuYkft+TtQPlhKCzAz
gsCq8U6R+SgUtSX7enGIS/FmCKeSLzZ1aYzX+sCIXEIiNPQEgRu+FFRRqSmNifxcrKWCzJ5pGyIY
7B37Vdkyb3EBu7QNgawMOgsij5Rww/cD5Adfs60NFiAlUBD6krbOtkhDpEnZudYCJWUAYkHeUBy/
whIhY0dqN5K6HJ1PD14Z8GuiwnTlFyf7gfGg6NO8cBGSUnQszy5u41YqVZMtvzgPmdpkd6zs+l2C
ucZLjooO9n+kJNH4pS9eAdja1PUG+2ZrKtCIRpQU+dWwrw0tpV13CMEFIR+0Euy2lvWbWw0aWV9i
tPtD9LaVW/3RkTg9lL1JTU1ZpPOZEU9J8kUIEoDLCdCaP1ztQJ8rRZF6wZTwRi3a1Yt9Pr8pamqb
1YHTxx94rJmsybbRJsAAI/GjBMJcB9k1WPxcRFgdKPrnNSB4gbbL+NqALgG1qh8MWJMzOSAeBVCq
4iAaA8QCiRRV2ulTEefHZR3RmfHWN4ZJbCxd9YhONjWITnQJyssGrMBm2ademmT4jytexyqOjZgF
kWgdPgFeJ931Zg9cWvq8nrsJvngRVK15UxKN4XbIrjvdfeNCfKmEKv6S2nfFKdazYIxe+qJd1G4M
L06hW3bzETNRtcEks4BTMCgUduLBDZMJWAjUcXPGCSTd+v4kpHOu6uxtlyGH4WeSIeiamUYpUQdh
OQzWZufPNhHi+fP0beaGV5PH74dE1cTaIZKxYF2+eFwsrd/D07a+giNLzfS60kkcilFJtrksDnmj
cWVMrEoRuQymYziwp2rXlx+sZC4mvNuPRnWIhjH9Ts5UY9kwV7UU9q513eo+Xy0+kobIC9NnNy9S
cYHZLIrzWlKQFS8cLSCOZ3PVqPXXaO+kg31mD6yKOtm6cUSlDphdS8IZ2E7HIWD91A13y1eGYmkS
g2Swsd3Vj17jBB01q5w7o0HgxWnlC34XSehmCD0YUBWIrn7RxEv5DnPPCfg4mMHu61ASifM5Zrqm
JX9MpNoOKK/MNzfsfN9CsAVAe8mmAFEuL96YUBGLOt33gLkFtdmCC1qAQY5zesRDYjWE+VvE6atY
IiQMsOC4YkRU65BLe05NAGhfQz3FCBVl2e8V9O5QsXhgbIT0OK/voz6kEuvKeZoxLilM4YRho3t3
k7ugqbPsYgZVQ5UY5pGydFmxGQx2+pv4NQXXYFWak1eIbrAKszQfwudwehR8Pl4WaM7xYALy9fjf
1zHkEWd4q69yssjxUu9pQ8P4GemwLoGc2JJyotkwPNbjUiL4vWo1HI++0yUboT1CqmoG0CpKv1n9
H2LxemyVoz0FqvEX2XJA/d96xZD9w1e5HGhd+/pxcib+6qO8b0KOgNgGR8LWwNp691dnkwdnHbco
I9AcT2bGfgwhP/7BbM656WMq/rAD+I9wkJC7CoaqW/3vk37wqs/fY+qpXb6hQ+F4JBgRjhfaKqtv
x2qqdijgQtNTS1rIsWy3w4AEj6d42nwaV3icX1FC1O3g5zs/DCD/HI8ogJp15PQquehCEOPhH9jz
6iWqpsnCEM2dvlTRxTsefp99oeGvbrq26SXr13Z4MtuXQrPLqDYwXcsPcMbG5JNebyHFm51itOS1
0jcylJYq4StLTvQGIon5+IaPcnEHQ/k1MmJTlo/z7aDohrBXet3atWaCBwgnDwXtDaWe7zO+RqBg
PhCkjahpi1KY01ZBEVAO0vGEFlXfuC3+z2ocuISpi5F1KLX2uy81i5sX3vgtykwVEwzq55eGykcQ
SdyBObHKH3yvAVavUMpQz5vPspf0XYli6+FEb/7hZFby0vIxhvj6ikyHVHINbsn+hEbZIA8i/hea
RaDrpk9uNNM77QeLlcasGkfGaanAgYAcFcm+7fJZucJ2pKr2ZMHrBMwCfYOD6l3tEZ5697IKf47x
2zkPErRy35iGOPqdykHCRTjsFN4j7KiifioXH7nnwkwGmI1r2RvudG10ueY8Pgc9grpt4wL6G/wH
TP8dT7veTes/Bdu8g2MdM0fK+e+Uh61EnEjcBbKbLVB4m/ifOfQD4Sm1756OmynpauFMeImSvRYr
Xa+wm5Z6EUGYl0wp+Ez9luaEXAqB5PjcrkRXJWGp5/PCxZYInV1Jt101wc9zdL7TjO03Yswv0qEa
XL4+xWI1nYh9UhMSJWKYAcGVH5E71x+qEK1OhwYhl/MEvzkhBNNgPXWWt9RuB3w/qnu4AebgH6lj
17vONYO2LRyiXpMgt9nQwzqsfmix3leVDGU1fnsWV0Uc8Z4uQHyrjgmo0MRfynoIJkk5ScBTCHyr
E4gmzA/mn6H1qxP3/v11WiLqs3Ga5H6MHqPs9TCdaE9i235Q2l1Xynepr3b2jGkI0ZOIQlW/M2IZ
Ai/JqPXTBcE9AJ0xEp/LkImtcOn5MfknMeyROrq/fx2Gay/PhbBuFevcwPOYRJCoIyJV5NK2YGAL
9ezoL19T28AyQ1SznwiEXuqrQqNCddgnAQLEZAhz9+FaxQKRFs1SC4EnImMLCT7+4jUEQvqeCd/G
pgQVFf1xqU4nRMaQiFFoSFsipVm124JjDChXjaFwREnExgwL66YsHQxXwRiRapV+ZGtY/6KdXb9t
ZPjj9v6TKYEXOU18A8z7nLNc35rHFWtix6yeOp6yk9F1sD7eJ7cF/G5jqQLc9kWgDvtPigt8WxpN
k2AJcwn4pmbsmZxQOITGto2DgqHXJmSu4PPGErHGVpzmKdAHPEIaOfVrXCPupGE/dGiMfRcB82xt
i7VM3O1Pjo5YZKGYseRbH+dzzhJbFYeJ0u4f/Q1Y8Olwd5PhtKyEGod0V9FsGBfU9DMVdVmUktyo
uvAjPmaioA5/uIp425dcpMX+LNLn2eHNwKYCwh3yomMSy6J+WnRHeulbiwyx8RztkyScl8a/Sje1
MXPQpahGsXKlHBC3K7Ye5HtHWzkp3OVSuSMz0itEXyVBeRwTgPN/m4sM/M06pUR4nw7Ysj8OkVQs
QiZFZFzvpS2rmhFQ49OfQAohCQ3LZFKkz5UFK9tVYFlPg9wRcX56mxte9o4XTl/1Q2huKo0XonGf
XYBZ57btgQzkYbwR000TQ+SEEHWxt45pooE98nLYuiOqCgMPUy6zUsfsESXcSgvmpeygogQrxXYf
RxLSFkmG+CBTGI0rtpvEQVaXRQJDNTD0IQVt2UBJN17JfQRLjrr+oLT4fn91k6xIGFfEnCXDkr+Q
WiIisv1Ze+pGxcFjwePT4XVcfLz6vs4J3k2QykDKCKZ6TWoeZ2mnrqRiq/tmy37QvLImUCrXnV7h
klOuX+ccm9pFgC4APbAW25D9n68UZCHAraCWYS/nQiUel3QON7XMu1qTLuin/oo0IODbM6WUws79
NRrirQUjGZsvdJuKI+geX9DIxi4nO90zX+wd7fj/CldvnUrNigEjWX4gb+nIh1sBHHopOjq38IZb
mMMJf6QSUZudLHJ7hmzOu1yJJfUmjr0jeCWK+P2ChxBdfeZDbHhXs+G+yYdjuH7oTF8gIwqXDR78
gFfkMgJw5iV3mx/LYPtbFq+3yO6ufisVX+5BUVUaQHvexrbcItdPSefqGHTLmJn7I+Zk4/8RNstX
NCTv04DeIw690cEIS3z/u4NJE5eLTf9mE4fk2/1fAISsIQKOB/ZGjutqol4LafHe0Z9Qke63j2kP
LY/f1f039VS0tC2F3FLrNSrnL2tiKtu0khwsPotD7odCnERi3Chly+OFNAlKsZr/JvJKqcmrJWKD
9LRqFVHV6n/7wqjN21eiv8FR3xTVafy6eK90wjgtAX8y27jQyHMNUXcctR9zW72M1Sz1G5eSkyO0
YUdIGhPoSm9uBhawrj4gek2GgugSD2ms9YMv8mgTHXEbPFPiCHLvMCGh0gsVnuneTxNYU8yLyhla
bOEbef3c2Qk4gLvSurdraNPfSpNFezfMkfr9JCf1W4M9vZf1X8QP1Hn0X6UivU2aMcvvWgIb+RXL
DiXhNDWNPVBotDBOjj/f+l1UCc5CsFsGKzMsq8zT4BSs4yj5MR+SlPe7EMljCbrW50cnXuJCiwpq
rV78ErU4fkT0KqVFlpzk2Dri4fPWJ+iGA8PLFcea8ggYY3JmIs8i+sC1Xe6aadz+6pbx1JjwJMqN
l5W39b0I3q3HqJhF+x0OIK1h8qHZJtY7MKNYDt3CmA0r7l3Vqbpj2ebWDllMh8cCi7TqO5F2lnxf
KUflXeD2nVAFnpikZ+VZ1Zb1FC1feiLKO9p63GRuscwmr2HBav1HTZ8sAGOzi9kM1iHGAV1oBD8g
zFB1V7p6Og8pbheZziLGJvnFHPCspGwZOt7KDExq7jWeV2c4NMMlxbIhzFq8qkygI4CR8W+K9R77
Wb/PzkTiE7qOYMKEziaK7JT/HUpr57ZssSYc8JEzRy3+oY9xufGqCFJMf9la/XNhAX0jbbqe0aaM
eb+ECcvypES8tZrhQUPLR22d2N0V3xKIiwrB24FkrkPaiuYN4SsKxOzZz2NPOROtzNdsyUNTKyyY
CPdOuEOGuaoIabwjEzHhU5eGI3rMtvbYsz5Rk/hfZHnvAtBTkgZB2k8rfIuF2IW/Pg0SAvDbWc2Y
Q2rjJFDm3OgWb1F/v0kuosORgImM2NzJehD6NJU/s84rnCLfNJ+roZeTkvpwPlHqo3+SBxvTBdEO
BjO4UG8LnVeAYfCxolauCZHdtPTtR5nf/fc58vkuMt1jkP3KcE2HwDztIJlkkUxCBciw8SiInbjP
UvKJpkjLF/FwQMs0BoWxvo683YTPQHe+v82CnUbDzI8ZOKevBmdw0+8aTtaokl/HtVv8/lWDc/qG
mAx2XfifLjkY3uek5wmp+/laYzaEbXDMdQty6XtlRdoGFEmtS9LOVw02mFfmxAx3SwtqdCK+7BMr
OATdRFVcu+7JOG1HWQhmFHOfzJJcniB5pRPxSBalJMl2Lt3pQO2Iy2l3fGB3s98ZHeL7yxJWxxDT
y8QnYP2CnV/WaIWL4kRT/SEihcvOiF25yUbx4jQVV4Cq6rPrdPUKxFTrOVWz9SyxHNINQZekDBjq
VK8GOGT+zYG2gYkOkH9hLcHX11sUtLW8lDVCEMmDbUwgl812AfT+fQ59fmOtXnHWSeNk8P+6XKOy
xEI5rcy0eDDQDIVUHKwwuPDvuxafSJJTG+haMVIfCpJONEf7hkn2/mu9/OnmyZeNYEZ9ZPDxH/TC
hl+D8BhK3Al82f7fOtSXzonuN7LKyI/sjmX+/UDU8XkN9Fk3m5w8mTeDbSmYa3k9/r/9AJ2GgY6p
hIAqpffjQ+AHg7KCf1Ezid6rwzh2n3jDqi/Sn64ERqEZthSd8So5Jcc+OlAdq4n/a7tHpCGEyMuk
ijncBhFEwsW4ExloEXhGvFheDqe5oL3pGJY9vI+E82fTAK9n+D54exLlx9SK++vu5cvb/Ystrz0j
JMfznC2lHmnQWLU+wz+y+RHgCbopITDqkUcVEqDevUOKlz60EnZ9os4nho1fHfVq3bwqvZTGkg6v
m7qwZwTkJZH0TUK6RMmP3Eb6z5thTLWWsG4+dw90LR+0n42PDOZ8hiC5ZGwWI7F9EGGHZx/oZ7jm
pkSISF8y2lN+MzAhb0iolIsYbo9n6KpMhRmtHKWUjjvrcwVO0KGtd/Un+ucbrUo/+oOnwmk6M+ul
wvx+ND/iS+EELzagCAFI+Y5h4b9Rag6eRoUAk25OncG+wWg+Injr2vsjxW3/GuEfyG9Fm+FJW5Pm
S4jf3rMoyA3x7xM2XdgEmkx6T2AoHiy8pzaDZKfnzdzKysZDuLFXE2CoyFF+kTgwlE382n0CLpLz
EQq39zeRrPbBdZGK0AzYWxJDyxqtkkKH8/YGQODIQNLQ34kixpsjnaSV5gQmqHhNdjKuTkTMZikg
hDoqmbuzvj+H24cYUNsaPgw4tGMOkzOzUSXcZ5t4M3xUYbt846Ce7TUFsunOcF6ZOvWoIbyLY0tq
9K7X51t8L32RN/Vfp6IuUZGZVRTkj/Am7nNKjaO7NbuZcruOoDKV6ppeiVClBdJdD1A+Tsih1aMl
u+7F1c2GVN7W6zBv4dQ6pgE7TJzSgrMAuiFPK7HyatIrhmkYrfONrn3WOtSOtkkueRzDpqHsHf7F
MvgSpwCBIexKIGeMpNfkibMq64LdbFc6+HKucX2SuNkxbfDJsao0x7igOJRXNgMAAZmHOrLp0dOw
9XvxcoCQm6rsYh/qA1DffTBy0PrpShzVhZWQaemIx1YUUAjBj0igvYe9OLbpEMtzAmgJSImGnjLi
gyWvfx4L4MCk2QrmHFmhf56BKdfAgFDMBc2QtZASmL/j45mprnxKnfRUN0ojPefR+e9jT11u+Qj9
iRDw6SyQVEG9e3oPGySSaRTqfUBbmtIbFesFdOVO36RSMPnxDKq3+G2xFun4fcgfLuoAEk3Yr1ob
oiFbdQXdhGB1tqt2QhORtiBJ4z0a8DtiHltZJfBqu1wPsm1myAGdP6Kz7DLTjSR/Xz7Iv0VGsKb0
A6A+iut8f6UVX5IGEnVW1gc297M8ykpx21Osswz1HD6GmlLt/k5wqkgr6py2gPD6d+MJY0jZibF7
3Dzil5z4SbGAXvr0BnuDy7Q/lI6CvG8WEtP0qGgXGR2expWkb9sfSYoaVYPB1C3hbjXDix810eQD
d5M0fkVF+9CXC2A0ocT+4f3lizENz9W2ptkrM3zWhsXjdnCN5QEnrv4RkcD1+73ECJ8OgbBM7WkG
T9j35PKLkKQKgEFOdtplZG2j3vpcR5fvFPO+cGIRccmdNpjHuwCK8PMWD/C6xjijw/s55bCbVY0s
DEtroB7m7AlgqaEDYHML/04t3yNJyRrTySuJ4LOP0zjN/8Dc6ofO8paLVkSZKTVJJbSLXBGkDsOq
9zr1FLZTSbLEs7pSt+I4QQMFAwqDNyC0E4EHz4lRj1mm0ZuzHm/kNtHbAtunMPtDNGwtv2TH6+l0
1Czvy+poFoTuqGfVKYYtwLU5ui2l3/z53qhx72MCBd2UaK5d18QNCnAbmoqqa+e12SoXgTibD9/f
dpD6PIN+jwRffflUU4EB5Oauxs7kJvqlbqcM2Sl54s/wVgcp2neX2rvvIIoUXUg5t7CgYiPTdbU4
mdKv5N2YNHvF/ByftV2pfSY7cRBiPw90FljLkNsl/0tJ14GqFoV7W9XolGIyxBtiOhpF2DM6ovUi
1h0pNQOPsaDXEn3NTxtcxjhvO6qzrzZrB67owI8oC+/VptwUs9uwq9fq/PtjPBpCF3WZD8wRI7NM
piOl7HOFG0USAI7mGtxlHujCgG4nK2w1GOGnyPiguh1WzZ6loOSUk9AI/l1c430Mkf87KiXpm/rx
sTMk5/wl8H4Oj2NsJ2Ew+LDBunfXwZtOAzqI/3Y4WZS1I/Q3cid9wi8F0ZIoiMQOtQkr1RXJ3aqg
OPXT/wep6//Xz9h1+9pJyuLKht4exR6D7XEyaAK6LdbFZXOFuTTIBjIZohPuwedXKmVDkwJoJfR8
knICHIOV4MGulKH8wXdT0Vjd2iuVxa7aOIn80n5dqbRiM/RvkMqRpHJ0pWurSOU2zWzlTWW3euJF
DFxnaImIHjQ6O+Y9/EnLffbme/858HyZYJM0mrRzAvfFpF7T1xP9aNrR9mCN9RpmnX9zGYltLQm7
hGbuDVKoYI9kFkYMr82wCnWDRTGRiKZ+fTYmnm2gjQdD9lMvV+dguML8QZM+2gyqGdBhmTx56phs
fkZQgcFIji+fa4mCsCZEHEpeVKpDkIOC8ap8WB17Mtpzt77dvnSVQUMXzK0RP6AzXWixGRRYnmYn
seZzGyvSCyDYY7h2xqWuQzjjdtIn7Ud9EvalMgqIZ7OsVZG3f8bkL49K97ivslfTZ//wqqDTIAcZ
+4nlAbNpDoCoJar9qTtXvpcelitYzhmM2x0iwt76QUTpYcbq/k0QhoDU2cyrkqJgC5wrJjipXDUq
YTUHJXCHBioC+ozL3lvE5Nnt5MAnZ78oBvoIYM9hXx+leNiaO5iCxUtYFbDN6dlPBvKvimyINMEB
JqSMfsY6UcB7iHDCZUbyIJwKAtn5o3jUrxKHtiBAiFUdH3ilNOrB4mBv1lc7GwQdnXZeiV1aZiiR
ue1zdbFX0WGydBxDlKdoalCeV9y/joc9M0+BFbFWzeikwHbqVtSasL4EvaFH1/oEJD8j/A/Ci4vR
i1QB12jfvUuuoeEzOkoDYTdXQKKiUb5Sh9d+RSy2+YbKpQ9A6Qf4NsRAtGzQuyBIzowQhO1Kcc0m
RuAbtSupvLorZqznf6aZwKX1OMiEaqa2VoFvNdP58J6ZAu7Stqx010iDIWZIwysyQecH0gurXqgA
86v5Qo00M38nrPPJ2rUZTw+uNXdXmLgWUSCOgzy8HX/CXtkxK2vGuCQCJcav9MIMBMADpzUIgKga
fuQ0cVzaMl/vmvlyyH+xfRK40wyt0q4e49bQQC4nAT+XZaST3zXTFhCz4RoUztDR4lMqEtiZ7VQc
Mt30YhLz+4lP1wqWBwFeG06B7klYxYC1XEc/2dRjITbHsa2Xa7ttom6bz2h5VcgLBKuLXDZT+6Ej
p482odqqV8wRffcUEaTU3XTUC/OKHIpJyfRAQ9HZQyC+DWiucKP9UeqUw8npjQ3hgUxjmR84x1uI
GOWpntNOca4FIadSEtNXXUxjvY8HUucgU+VqzuHO/aCEaVDMRf4BCo4L7nXm0BO7WpQRI3WpYIbJ
HjhYOxPh+clHIQMUWv0O4wYVXY5JDrlkeF2Yvwg5P9yryvIHsTM4FHosJtccDaFSv7vfwkzieZS9
3u05dWlwd5O1xrm2oALDf4SJPynjwM2T55Tn0iDRdpJncWqZRyTw7zwKAUy7dplpfVFubk+scahr
74GdrAmMYSy/gHE9duTZKX6tvJB6L9fckAClydAtfj6eQHFVFiZPqDH5i8/sHpFA4fcXvSAWDDy/
yGnxhBbRBTt79eTfekcrTI+CikZDqHO+7KPif5ebiTB61b4H57CFEe8hbUbUJRzm4r7BwVHPirB0
7Yu3zHNkIYDlE9DVndPBWCRAk2V/LF/8Wt24hMkk8piujH2GvBnPKwt/Dot5612cg2qLNSO4/KxO
SbSTpBqvU6OCHSc08qO+7FlhBZfb4O1fyuQuwciHtdG5tvZIGoHuxq5oCa19u3qx4JiSKqv8d3dt
JSOxeMO95CDYzYukT5iy7mjNk0cbn5shufrrwU0i8FtjHGhD1CNpSbpSguzQ1Jn8QN3uNE6PAM2Z
myM8qsnk+d03NhO8EAbBvA8p+RZTPc7PNpeuVVcrqvibfelrgBR6uOEVsPE8PKgz8bPISA8p8CN4
w9v5jR9PcvU/wwy3S8qNumFVyTg4WtKgWxBRy5ucm4oa7HWYFyK6PDG7ZxNBL15mtHJdtd1IxH0X
B3IGsazaTDxFmiX0jzmayu+BiB0VDzSe0clqALl0yCyHMCSXZkpabCTQD2EVO6Fh++472TVvL9PU
Kctgspo7FFsiA8MeD+soqngw52Uk5NG6zsTNVksQYdJkRFdAer/rdxBACsJh89AhZJjcGYTCa07d
/1aOxcAs/Oz/GWWZiyE5MDEiV4TxUmi4x/ea6Zha6v7MRZXdZjoONb5jOducwWSNddYF7oXNiaF6
8w7vf9WLY/mE7AiiSXVTzzaxYKgbRgQGyYemWz/fKbjIkYs0rj0HFovn+q45bXa7Er9yTCOgnM1w
Hk2SOnh73gw9qr4w5zH7SDd8gZ3yXIjnBqKow6Gr+YAQ+vTZ6lpPT7sAoxlUAMNtVW0dIXbm9dQp
BTtHdPnnggF5SznrKZmMtgBs5nMMTMz6D2ocCquQfUhZj2Rvfvd+/BG+Nk0IKiwRe1zecxrDXsxY
+DxHMPZ4aRGXboQ9Xsk/JyCYuJLyCvo85XFik4LoaqQWqXqIxMzNI8yX1ABZpzR66l393eiEUZTq
noA8u1bwUqy0Z5XZJ5geyfzn2DrHjlMEWbx3T/h+un2uMgXCXvNG1HO29qX9EefAOwOspmgTFT4e
4hH+xHw2N65UOy6nTMSco87P3RzO4sX1b8Iop/bo449m03P1I83STu1GuGgLztr6duiApXJjRs5c
Owhr3t2A9E4KnzOmgESvH8qJ9ZS+9owinaDeNgrmZKAzEyaMGKyq8HTn2+QCx5kR7ANMMQvelb45
ezbZrnzPfVMPPaMsMLYkhYBwdqymKxOY7fEVQ7fmsZ006BdRgT+8WGjEnvggARRwyWEvftGTTcXS
gwVqpr1XwFGKgN0tQ9q6t0pkFppF8kGx+eDjUvg+fy6rNhYN2nDgHohJiP+YbMUeRLCYVOilL6qr
wS8ct67+jYoN77qmKsJWuVJNoIthCXzBdNjd72peSRPinRxiSjog5VnV4j2F/qWb4yGaWK7uzaQr
12MSEJsLoKfDv/IRyGh05frdZMip/7Bjv5njzV2DRFTsrxop1pt/lbMFSB6go2cSeRpsPuNjRzeW
1K4oF607X/PM3LT0Hwiic9oWvap23mqeAWCZwEVyu0saCUgCUan6rEe8Lx0SmEeSaHRihMPVfC/z
+Wg8m4oU4f/im0QIupKkiOODOQL9wDrZEz49cHNYHGnqaIK3FYTN1n1SyhmY//IQX6f/YXfumbLx
+xk4B+xgDvWbTUT4gfc0FqpV6heyXZYPAhdOSEjmXC8DpWr5MZC0KfgFbQSGUoMQoKkR4zA80YC9
CVgqDVS5i82b8Le4JIYIn3D9mrnSwnwLqX6R+yegAlMkgctDNuGRc5COf9JrAjBCYzSJ8hd5VuvV
dhM32dgMonJjUTadBZBXJUoXtFlVQRIo3hqJs2mWFf1fBBA91WneLRLZZdP6ABhCrZpN+B29C6oJ
LJfmpPZkmqSAV1uCl2yeK4UY1Blv7Osz3zn19bWIghoBp+06UVXvyQe2v+UdcL80F4EFtYQD9Th4
Yri6hTk9LFQScrsmczmPU7IeadKl9Hz7ypZLUJCBguQCkePBd+qluqfJfXz5pCFpCaAlWN2KdM6D
FTKQThMwNgjMQ1NQQtdQfvKbLTDVBqsmJNIfkt9o+lrSVMjCPxqURDlv9aOY+NEoKNUJ+D16qgml
6pbMmaK6dHoZjQIoTVx3FWqXMfGyxv3YrmIWaoS4m3ueVCvXj5y+S1FlRaatwL7xg65YVHpnnbdL
kSbloMw+gEcOCSIUKEGIMHO9DvnRozaRjKLmUoZvUifwFDM0LPoDeDrgfaN6hoSCYPPIxvlH5PAI
nKTTx35TNfg+U8xnXv/qbJjl89vVSeef9IYXf86prRq3cDfQTSxI4H8lPjkOa9YI7NmqN8xcGjiB
jpk9OMSLhv2cGMgUg+hQUyKrxDnEQtCX2UwE5qtgDqr6Cej8fc+tcRIhF1Ux8S/4cUa3v9Of4vdL
ku9GaM+RYKL2XDU6g5C9lFPlORs55ZVg6aR0q833/ZEZSh/DTh088QmiMG4uWywrJWuxF6oGlYXw
DOmwwtx6/uWsXSosDAkzzKHWmopgDVFTs9BnvuQqJyrqlWGmIrR5CH15CsIHpCiuWS1LQ6EXzGHJ
kWDP++Y/uNVjNTiHRqTt7AE9tO/h2Ge6Ho4QK2FT4uzPMw0J/DPOsSyDjNEvDlqImGNmS0KdIsSJ
7wFdHLo6WKKyvzLO6Eve/io1+V8kh+DVNoAKEVqpMpkqi/hKnZm8my0ETGy15oPel2gzR5MAUX5U
YpUgfTj7YmmmXBxHJz4Io62tiZGXk8LBf3gT0Ov+JAxnfsGspzFr8Ov9zjey50aTly560SLKcTey
G0FRKIZXjpBl+RBfqlJyWbvyGV7ZTu4wNph9BTWNmeSz5in5OD5tOVW756k3cJndXpRHdaX9HKL5
PXiTjGbQgimBosN2cmj1t0aXWjINq0Gq+t8eoee+K3X0jMqebEflh1WqZmMoGvJmcWWRsHW/xi1z
vtBP1fuhYS69NEgK9t0kr/n/rjK5dMudOzaUGlYjZqau2g53OnG730w24MsrVjJWdDgqmpzBiN8l
JmytdhHrarr8zbjxDqMzXy3gQgfXIvPdqt67KFox0TA/lgvWDebpPES7NivkV4WxaNtCxLQPMCIy
EQGtV2Zid7uoNXBvbiyglOneFytfpfgZsM5TS/5hfwlyz+N1X6J4R4YJhVCIKQ/CSuz3Gb4pawrG
Vto2gZCi0eDt5XA8jUqrpHz/iDtbmeozU0AUUPhQyRK4Fk/XYzdCa0D+E3ppJnIZgg1qSXOCR1qU
a80GMNbN1YW1GQDC5W87Rn1hKSIz2ZT/X4w50cbv+646DHvXrJkyHSpVM8rv0ftHLoEVPeRRC/rL
rp+lJz9Fpd0Px6B+uWk74dxea6coXlYY4JUA70VpiDPkZDDt8YZn9ZMeM+HflFM3id8whD/JaCFB
IY8lpEdAo/mdx2pFWbuk74SPRXV/IC6eVdhFXPJLBbTndqgL8w0I5dX6nZZR3jgduG9W5kcn51ak
2GM62mVqiYi3eykazaZxIAaelZVXJn+ktnGTgQu2ersUePKw9/2qQCEBc7BwZVoGltD2uREqhdri
h69LPPRtJkhGYSgEMSlkJVGbEuKcOKk7psDY8kEZqdhTnMpBsNCVOoi4/Q0prYPXwGWaXcp1HAvx
F3xDmrfsvRj31Jd5091z1am+wZ+h7zLBscyFmkgLrbJ/BGm+jM+LkKZ/vpGxKSUrLFZWj8QDtoWE
VHocuMlHlFfaHZZqbHMbwazmmWv/pNnMv/jqVX33daz5Mnm2zfr3iH14tpUxQT60NKtD1WRuLNGI
UyBuPKfBUlRe7MOPCb2WB+1kUV0HPElgDtDi4eK6KBPWWa5p0erfMu0ddfjGWUx3Ql5hhKt+w1Id
KvDc3M9/1N1r9ZkP9Ga5LbKV4W4Erq08oXNJe6qFI6yTGtnxd1ueWX/8yaMzfWyXPyZKKJnH6/gx
xG/4mJpPuG044kXVD9N/PezvdT18Saq0yTkhTQbbvl1+Bs1AI/gU2uQbPOBmRh1csPBSzvDe6kOr
ZpKOcApTAmAkN3iiNnGCFkXVEVHNhD2jJYg1Se9RZkEFQFseXJ9t+fVg7GVpNns1ti5/GW5TDrFh
7ging59pc574FkVMT1iGJ/OLdsF0ihVJYnxU2PqYw52qbasGjEvJz3sNrhQ/Vw3hjq/TwR9uVuGU
ss6GTmajjCkxts74M5M9eAP4BfigyC5Uec5oK5m0cytg9i0l2GPxMq/gqhmwknQfEHbALvF6Ht1c
11RHHfpydkAdnsBJHVe3ZudIlvTQmQC88b66c/nJ/rHhIHbjd6+KcWZABBgyefnE3SOw4lB4pwkA
eojA6SFy/kyfROB2KhPoTEnVrBk0ueUJBJi4erFpd6SNaHKBJwBLDxqyx51HZmjf0fQDOq4dm7sn
bHuTYid7hODd445VHjcbTuXkxTQ2ndlMolbGuI7QDRWXOaAKOp/ayY+glr8BsIZyW0hDpBFB790p
ugM/Ehrj5DWjelCHWJV2WGwpHqLBo04jCTy1MS2JM4eQ8j5EmGoKDVYsDxKMQOkDuPZNP2sTaMQH
lcZsGUmyieDjErubFc0vJitThZSsJePYyRdNE1ja8GbsS/tuAgL1a54Sada3rCzSiSn01hMi1cRp
2qaeabpi3LLtHGnNtVwzp0MKHFqjzaElzGFgEHi+hyPNCv1Iu+lWX5c8FGE8+j+tRk0xJG9++Maj
bo+/U8eYlJYl1dJmK3m1uObXjoF/BCZbo5seNbIWOCtB73SZSuEIv5bYnDFd7GmZ8vH9VPCGSl50
g9c6MnGVYbgcp4BkHAm7Fo8KVpGUdogzYORgI4kRC+8Au+0mJHY1rOjDicxdf11Tt2A7xKm24ljK
WKfuRSB1rEYgT62bXR5IqviMGEsZgKFy42ju73kZwsQR7cdhJrqlYGKLKWuuA3ePYIgHZbnl9Xui
6WX2uJOXI01lZ9bm1p3D3yjgnXgk851FEyo0L6R/hRBN+Ayhonfw4d6jdDrA6qDj9nd11KaKG2Mr
qNxfHXTjrn+9PhwN46u7htc/Tw1renAX3zE+um1gJW+ELC/knjCSR9GeNJIX94zJ1gb1Tqghx5CC
LKR6yqFxcxOdZ/YbRxyIuSiyVafq0cOaq5Z9c0KbnKAC2xEksQ4y5Y+XVjeHouZ/7Ud12eljrr1P
pYmXXHSa9SlJZM6sW8IUAL8cGkDJOmRR8s/9c40dz3kjcu9wyzKVdomeuNzZ8Ytz14pkerxfOmaL
f7j5OC71O7WgSCunqYXZD3VCOsyA/6/UmbUljgVRrD6LOjKDw+WJJIgKXRuzCo9qAwm1Jyi8RXSj
+kbVwkFXXEkatBbv2jepIUBlDaNkiMtZoqEmeBy+T/2TDqeknlfb+RhswBR/ahWRXU5SjX8N4AVW
4MvnG+T7jFuYuGekAzYNvMvkothCQxtk3jqi+CHm2D5eZ7k12xqJoSVPSzx27fBCf4tIn51tQg1I
28O2lDC0DwSVdcmgWpS++pIIGd/IHKIvHqFkHIM3HAIVsR5rrx8jFShRE1pgUdu66KDIqgt7TNyi
cTp9WEdv1TA//54mX6PKC+XlwY+lXsBrBX4v/P9SOqau1zRTlQvXzOxIIQ46akUhc7Ov1fBdunOe
ut6JOCv1fntlZdvVoSN6fg6UvBZfkrWp87oS+uA5y80dwc2DiQe8FnrtXJZBehGfrSdk6zDXJ2zd
IzcnQXjNGAnEmJ6k4FclDCCdQ6qNEPOTuKHzZeE+/hC4Jj2Nw4sYeTxidqXnniui/jc81EEiTq7M
2/WsbyZTeLwCfDeMM3woweTYx741XQLRYrmHFW37vLXPDg/5EsPI1KQqJwhxnXtwY52Gi8p3vBsI
Jx6xAyjV8NR2A5T6Pkw+NgM8yY+3go0zvJ0VXJUoTIJdrDinWfYi8j6JtT132iUVaLP9mnu1fDk4
jxKqCJQ9aPcEd/t/gLhSMA8z8dLaeawcrsxyjB8X3P0JObSa+0rsTMmDpp2UcMxwGIfbXcMAtdY0
j7NhZfwhZXjhX4g1n4DzTJhiml+VyduWdop5Aen51VcuhOb/EJ7cthDde+0Yx/6VK9j+vdHzswsN
WD6yIkWL40Tge55cZiMB2LggcW+uCX8VfajmRkZWQcyXFap0BuRA2NENNo+fTu6tGp6izdHLMnQb
NBOMGdgQdaRnTG9qFjkcJaN6Q/hJkIM0FQAQuwzomguBxj3NvF1hfeTjHxiKhbSNKE8AWpgAbviF
E9hHRp0dKxZrNh7Rb5J7gVSDikAnz2bzGkKbfexUxxHiw06BzaiO6EpwBTFPT4+IVO5cr70ez+WT
PwilTqZaDOib4IRJCOXsgwWebXYd9Pimnm/FkGyeCWEUCXZxxuitSt06faOsF6euYWzeF9s5Uacl
38EBZVsobhEpF8Yys+LMud6ejhcVjfaYUi+1+sdAfFv/IGVklCZGbVj6z+15cIsTW+hrZYNlFbyq
WIntex6a1lxVYh866372oTHwtk0R/1kcCr9sfMyXf7ys1jA9hr44PEIySN0zif9sGJzDlHxzLukQ
dvOBMwTnOjZVqTju58I853oPNng1aFXT9/R/VTs+S324xAST713M/1hiTeL9ncyYI0g6906pWzgc
NS/mL6jfd1P+VmyMoWYBldxXqI+PypMRedOCY9vubqtweydxNVY9Cw+J/RaO0jEb+ENpR2Fn2j14
lO67hwnbH3r/S/wEUNAcAlkMf6Jk7shxxSjpsTiUo1VmP/Z26bucDBxK7ljJ1J7zYwU+UBcCaQQK
EI/+PrQo8wr+7csES161CByVjLvCHAgll9lpODX+1jcutFdzO/gR3kiODCi1sspuzC1YKmxn1H81
ROZv2vxfgyZbVlcUJR+qn0DIOuLKiXryr5/y74otssMIMcsjvCTNqlIMHRlXRv5BI1YW8LNLd7cz
LJCHOH8+IW+R7AkRhlnIum2/4N4DehijNGa6TEjN2lGCSTxHDVF/g4yu9BGp9cTQvCMEHE8l5jE8
zGWq4REVBl+N0W+J78P1MKXUM5oEhI/Zl7AtNA8zZ8tSzu6/RWcJcFunuc3t2lU9YYmblOQ2zWpz
BRYrU9fioWjuKVC2JcoVXdEjY2QSPURutvb6yaxtMrnP1grRGx1dC1ubgGZNsbHA71te6Gu8s2uR
ahy0ZLrJ+rOcq8SWmtO+Ch592s6nxESeubOUeNFC6YkGp+yEV7+rvcJoRsuttxDnNIVIvp1ML/zd
iOdq+4WuckylWQ6hzE8rnynFG4jZ93r9aUn/CudJr50CgeP5RWGmYqqp2P/NhHNyW/eBYUhJ3ZCV
G6760gGG3quzvtNOHY1G60bzKgY/vm+nJ1N1De5Y0/HTWwjL77TsixYTxyE7InxAYSSjH9r7f/cR
ODGIHZd1rDrv27u9H9/w6RY9Em9sm/7xpXVaIv++XqtzX53TtE+tSWFx8qA8O/H3BF45YJc0GuW/
WRvOukELpvavYRM3UTp7D3cc05Ga37JWwK+W4SVjLX49QHE79miehW818eIifG2cYORXZ2PknMTT
yraaT23dZdTMiswbF36LdBtzXd9PKdXbeFnTm9lXPv8j+ZI89o2jHWMwCi+Z4Jdvmdo+rFskx2d1
xAl4p8tnr/01qaRn2gJ5BEdRU9XdTder76+MuIxHKblzJ8sOJifhZQDSh8lhwdSGUxETUa7eF5Hr
nJQOsWpCLXgxJq5lBNdvaecKV0cY2huhcUBepS3urnf9+mCBPqPu2Xddnxh54jaxCvJfqRBI2Mlp
dQcc6Pmn1lV/BmJlFMAwOEPMzCygNKLX/f1W6Ef/ZCasUsCBWzga0gGZCikzT0fkMNZAlPwTawPV
o567y7P8SCEmwg1luKYu+5tjH0Bjgsd16BsPEPbEiJc0kBMClYQEhP7nKRdXALzX5mfQL3WjBqHd
kA2suI/hSC8wMEdDwRyZ0vLHeKPCWhk7H1ElsY2Mho5L6bXXDZj7zFdzePhenoMT38vApNtAMNsw
x4wnScZtoqpE52JELvtqY5WPLky6pDdvhWK7i3Rbaa6qvJtc7jzEEZt8KozyRRdsy2nEFDpcTQLR
CKKl7ABlwjDE5quDTn1oRO8uiWOeHbLLASrP/ItBR34gjd6VMiPAsKNCz71T+cEoOl+Eu5eUTskc
8vxijNkTcjCX+PbRr/WAQODpFwMZcMNDthKT2uM2j8ZIchGq2/524bxbskfQ6i5wpBVLu/o8wuQA
x/BVOwVmJK3GAT+ZgrGqiHnX+AK8iRi42/EHuB0QjE5g0y7IKkNEsqdPQs3rRUbFCi0W7Q78UevZ
dsH+XDYZjn6pc6AV60ejIMGOOzYD3VJHBp8Aq60qn0LQjizfe6KNLj4PM//6SfAXwKhnvWyFJInj
8TzHLNU1g4KN21kRL79jRIFn/yPvFJVdp/WWyVVOhC7dKN4JUA5+SWG1tjpkxQHTa4n2FxHwVRMx
X93UlorThZnEq76IPNVLbt1i33IYp8++DkSpPNCnrmr+tRuCYTrp9r6tia5yo0cCydASMIdcPvtb
d9Aivj2SUGhnwByDyTgpaMl9KYnQOBtrCY+kqET5GEhsdbu6Jm252N6Epc1L/6Sr+5KgVyxYAdCX
nWRsY7xj6S5tjQ0LafPOYczMsMIpAXeBBK6iCB0uDkFAT/g9bbMFV/GyXvrC3dW78IeUxwFgVlyu
SRMdLFBGi1HE4/Y2d8Bd8Nf0MXmTwzNaNC5C2tdP/M2lzc3LDxYJ/exdZvfuDF8kFgbxMnQU0R3P
Wuy9OnavdZhsgFQsY5Z18/Spt0VzGx+rJGhJ+6laWJmF8xn+5RWvCRdNgxVrrgcDSHaJJ+v6LPAs
EsmCC5/hmzrNTHlu7b5ZXq6pdpoj0MdafWYrPLf59VyeSB2H7yYx1SAOB3USEtUoaY1ETYTeTvdt
8duyGAfXZt55xnT3jmW3yVUK8nWdEPxuJLsIx1MapzGV/4StbVhLmHaPeuOLatUnHlpqlr3omx+C
mM1CkBd4AImTw+RMc6Fin07qktau8A6KGAAqt3ozOpvKMp15+aq1an6aPHrvTpKzcYV/p6+k7hQz
oUl9Z4mfzNxKaJVrLVPjIz9J7dsN2Euv7R8j8VwxAGJ+3iXNwYA2BTww4WW9Mpqh1tT0XeAaj2QH
o1OGGZlHJqmM7VB/oQ+BuljvjilggjL2A5sPiZf4S8NpO5nLhnKhgdktfA+pR1K2qCtl9tGwvEfJ
54S03BIYMav6k2o5bnApD1SD+q+CQ/+CwFRcOZLuTjX6DLKHqGRoJ+DJ0v+bx7uMiu7iAsmvQGcT
xGXfwIhgNwPbWBarfgA/rKSPh1QVUtk3xQsv+J4kdPLrFMy4URSNvTS7nmYmN9zGdYlNvOFc0HUJ
8dHygbog4UAjN2IQCHx7mlmc/N3HHFFAXshX8ZKzHzge1VTmSDSN+i5trngyAsaCDrqpnuO4BOW9
6NWFuPSvgVZhgVL/l+IKjfzrDuusU+OmOW2JS/QvQYpiw2eKCx/JQAe4pOovFeaoG5SBrDyzu6Gr
4q4b3qa4eR5wzWZ0cJzK8rzEKT3TxOCOrE8v/isRftu4h++OJ3eAbi1wJQVhm/esq/3/NRGNE4I+
ZQ5/aoWkiAt3iT077gIUuu8NZgvt7LtpHxFTXDyG6++zwzQ7YvdvFbVf2JneoCRivj8Va9m6XqA5
bEk+5+NIU9syxMekvQm6o2q25p9petbD6pBAGHxBDrCASss5iNhpAWk9UTBfp9/dF2bWcWkPjhoS
bEL4yChk8Zkm4SX5EO+OpTVY44bD88KPF+CdOGR1JFu3q/+7zz5FCjJ2zVlUawb17uQa8mNQHCzY
cb/iH7xtvrXoi6YZxjzFzQjoVqLaObdz/p9Y1t0xrBvtPI2ny4L9cK9QjFRyrcwDve+PFJNIGbGL
84lOSGemH/jdzVR9OGTAH2d3fW48dxQ4HZxYbvO8MBAwcMJ5FXv/Jy8upfPAhlnUdRwGRY/NVcxI
J5cTeq775jHYMamfviP5VjQHPOtClmfIb/IPyZD+zKkZVc8PdI+u9Fdtak3UJP+EQRsyEVvQhQ19
cFiYMdcDiBuLtlangq6WlyQe5GPehM5OMILEA08Wq36TKzzmqaKPiE24JNP9qSl00POokKAH3X7o
o5aO5UBRaD/EMJbY/cW/dnBcqfiCFr6foi6HmIb13bEVi07nI1iUvIxT05daNYpZwSti9HBpj91E
pbZDt/Y56Qy6o/w8G3X2KMVJAkjTmKan7se/X2OFsr5mtqEPsjNwhCkncCWXkuEgBSNOX5HwdW8u
mwA35LD7WionxXLJ+3LsJP3Ftj7jhGFM+zZBpU5pE90JfxAncAJ2kCCKz/hc55uIjWsF6kVkt/bS
c6PpXIh31IxovfJYjhz5cgOwzEy1fFi5Okl24xGzpkCcW5nX+jH9HyrnW3Z6jSfx0XJCsN0xvOd2
xp1x1NpDRJ6z0lj/LmM927ig/3Ey4kK3Y2YBMCYExURvg2KzQT3oiE4zEUGkkNdfh3XdqWwDjBsW
FKCYZLoKwtJgVwK3wni3oQdSPA9NQObMxlF4QD0h8cpI6DnyVAR+TloL2gckJo5NKIN1VSnL0bmE
KknPo9sO0qD9R/vmxUg9xXHP3IndluwOKgyJd/MHNHZ/8XIEEf1KtTjVuMq8zjsalhSlaRlqEyx5
RZl5mIvsu3iVfpsHAlUxE22xCHrs8zJgtt5QJzcG6I35loX3CsOkDTqQ8aHqVgJI4T0LYCDBPxjj
DTkUenAyXUXJ4HBDgXb9K7V7alYdrMtpba9qIkALEGrmxeIUoOc0wYUB+A9dRJ29lnPgOdof/CxW
RysWnxKA6Q9E4UWDCpz8KG7oAykZU/tHdo60Jzhx1+vOqDWUV3zd+7SzoAQ4piox+/1NHtoWPZFP
bBJMwotFJMy3HWUOTiBTUOkMvYy6WKj3siZlKeN6WTkpyg932c2hOvq63lpJq9IjFK7j9YSVuFfj
sbzPbA/ZUDf/0VyFL8xAZbmkyMaaBBJLBKmwIkVSXqtrGVFsUF2O7MzxPLqu1+tq5y/9wBawbIBN
l9A+2akn6bl5OskTXzdd2YhNm8flZ0ZHC67+9/1Mitq3cS9KrbRR1uWSy4netPpa1L7nuNK13hAt
cxqyzj8jbz7JPqETLy+JKHsyREhap2MOrjMHTkHRNeitGvocQDopHq2OZ51wDA6YLsFJ0uL3cCcB
gARvOJIOwU3iMOemotGImHO4Z1YUv0clLDKkcM/+1Eueh3QfjTAupRImSrrLoG+aXAB+x8cJD1FW
sSow4ybmeqi+0I0IXvwwo5xUVbMLXNIV+1tRVUtsig00qMqxacy5zIRZQ4uVkpb7PXJyMMSUygRV
d/8vrGPae4HO3iEo4he3U6m80S16fRUgqw9HeJpmg1UKP5iAphWg1g9bejJjHNXODM2Q/igtV7J/
usveRvUX21+U+puGvvBEfxjir/yDhykKfyctbBcpVeG2bklrWZfz00u7RoHfz2P3i67n535fmYyc
bs4c6W0OjAD3o2FUaiQpp0f52OySkhN3Jiq74CSC/N9c1KmNzxa9jY937jjJclwKnLNNVMW4bHcG
tTxgnzCQ+BZ1ZFViri8H8NWgsyfNk0fvtXmsnsGG+9EkQ5ZvZxn6NeXJsEHSn17To1IOQsFb8OmT
ocbBTTTRiF9Qj1hovSwc3/mW7c7KuNRM86ZRQORVC/Pna5ROCLxcQlz57LMc8JDlp3tpqhY9iN04
g3Rc0hu1GE8uS46wkkm8aQkE/iw2ZfGeA+o0RXwLU0GuMPP7m5w+5QLdEsfiF5Ceq8sJKyk5o2/O
xnDzcv3uVBmnhMpWSC+VZzmNbCr/2AdWTpdZjlOV9WY/eAf4ooy5MuHXlCAQt85eYi6MG3aoSi4K
5mnNQFDYKkTT6Io4HBoPXRi+7vQrh/cBMJ/Rf5dIQrkXAyKFxSas0pMfakE4Ldyx5eDa/9N4DwzL
NRWD67Ks17ojhNd+3EV9zkKAWho/fmZ+8QJoENLsUww1KGW8aQL5rKtoPbZpoiPOXK1SHK+yo78D
zcsY7wxVZ9yXh3vfEd5dgeMc7jsFzXodFU7MZdxCTntyYkq4vUB6MPsUrEOUjvGjN6MCaQJ7qYBD
j83LQiiWaiBJ+rnVpjC3oXR417hIjnrXFCYsTB7XGRxGfoqn9YeilIUcN6uom7dmqWMxSH/1qL5l
f9CDUzmMnLnADMfNH26puu09RGbsL0A9RBNTSkRMdxRVcBtuDzRJQn4Rw/LdXJ8/n6+L24ci9/SH
1Cq+NshHmd3Yppq5BUijpB1qCzWC+PVGJdcRYkkMUlEDDUNLUNUpyfRrizgvKzaBaqQ878uuBYX+
GyYKvAezy8J/Y+J+R/UkUoKracYTP8zJpOdopba+aFDjZkdPJl0A6Hz+mu9ScX8nbOOvqYY3zVBM
JATzh+tc0yJ08Zm3dvdawyLtPJJJ+jIXrDtXC6/PPUh+ZcytAlZ31Uh80sYPRfDMwZmhyUx87VAm
RGa1R3tOY5jGVOawjws+55HtwYbosd12QHNslJLh4rs3YDuxsSIoPf1HN3CjZwGFCusLBLVoQ0qL
9PwH5p4x1DqXLidD4W+uroS5XnDmugJYcMrfLtohKHlpiJ3nVzYwMj5V8VT16mFSccaJlFsXWMLh
0vDOyBMx8lzYZt5mEu7akAGDeA5COkkxA5YlIClrga2GVJyws126ZA/2bzgHiAtdPnpXoVGXKBr2
2SiuDnah2eTXFbfqz5JnYWlkaFbPDhDfo3gkcsPD0Fe2SUW+1wh3QtAXAqtwUSeiMNN8IO7a0CcG
xAoIJA5uMwWuNh4TCl+hDMI3Jjqlei30XG4QVbStXGkEooPlvqu9rxEybE+i33pupwlZJ46uvMsB
LEvL+Tua0lp1OziAEpeO0RhT/ZgVKouKnKh9icvkVokPDzxU8b4UYYHKzLkQFVMWCkSHdt3T/mRq
zp8P4ubCE/Z5rKF2NcJ7aQ5WPWIe9/o2b3Fx7EJuT2O3btq+43BiTtP19bsKiG5oaZDbwAQ0Ds6t
JKJHqZWW/Upe2ZIqHoylhsHFWLqfzfV6JLY2jaC3WdLdpb72InNEER042DsLBOqm3tS4cbAlzfuU
Fs8JIURrB52KiHNd31TN4w1bPNy+HhWDpDajeUZrAFBTtC8g6+qXduTu5of8fr+x40myWXEq0GKR
vvlNA7LxNnow9MKvKd2N9Y+P+0WkgSMy+sSFgyoP5YiLxRNZIdVS7MY/L+Fyvep0SM9HVOGvCpHN
JX8YPWKet4aw6V3EEqvNiQwv8pY3gjX0Oit0y8Z+sh7Ytfyl7o50VNMcytJPAbJfez5NZyGnFRaI
R3uICqijumjEmeP/hPJCivGIwE93HYm1wVaVEgdTVLvmCCHXL/FR5csV1QejJrVpne27aL7FLXKC
j5cXQiXD8VDjhwyhdDlHE/0I6RljfGZKrASH3DHdfTuLmjTV8MLgTbaexbTBP+TYzIk9cHbZbxGP
eB7agAjO+WEkYJiQPU6Uun3YRBl8OtU6Tw9dzHRbVIiqc4m/B63HelJQ5fyEP94LDqwP4GVIsGvp
AI9EoWqTig8c9HW1aqek1cjD4y1Ni6KxOx4fnRQix4XYu0f4nIMpE0eheT9eo0H3TR2DHTmLI6GX
e04K+hGKSDdTEDuG7ghVfI/l4j16KbYC+qm9MaCL6bX1jBHnXyHSKR3hpZOvRyqvPxMKO6wy7OMp
ccHYxI+4+HMUvevkYCk19eBsJSkXZh9GLLbtzjYKOxwABTRcDk1bnmpLKgbhXWXV/axDbrNrXCAf
RTpw/wF/0uiJBqIDSQ5xvjuSeKQfefV0gHQaTvncX6rr1HW3IOf2M3s+BKCM/pWeTxb5jfFmTWRt
obRcv66PdyJBgbvN3pgSNcxPakYoghEcAv5uP5mEfQ1cWBskIo1QqSKJek2QgqXhW6nIljEc4fyl
eslxmZSue5ZwJ0iFuQkwY45+4ta+IvJgYJyEQ3V9VW8F57HIug6Yb6cFYna53mroB6F3Md+xc8qX
JeYxRO87IuKdbQIasaM/Tg2XYIDuafDIRFeiHpp90pGnMperDwhb2zOGznusH0o6UZDKVeFC9j4g
23puFHpLJUQydQi0VJ6E1lRKBEbH6VSi3mQDpR6dYJERJHPralx/KFxrsEBp7wlj9zNqvIAQ/NgX
Ui7RPee2WNwi4ba+L1CQcmnUWrGsB9NqiHP40fovkFdKm75jXeysGiyrPVTFi3zlJZh5fZ6SLm2q
eGqUeIsJLy8D31Wm9YyK+MtnhzFtF9j2YA6cEkIjTQF21Idqu9wfSCpxnq+zqRAzHYMqKKwBlYWt
bvxAQ6YDnmwqlPOJeAXspUIZLh7dHQ6YgaIQ7RYLbvUW7qzMlGqorpSZNOdW006CXX+SZKknL59p
ip91cP6MN5mhPDCLsIBl1C+glXy2pti+Np5IVpxyggd9ZrGaHsL508pqQtgOu0l8LW8XsYlYnJSs
eeCFrV30IddGlMfyfnb3YEBJjOUmwB5NDEgfJMWuG73LakSJWJaoBcmjMex1OTFWe3MZjaii4GvM
9z23YGYMwjUXDvsLRbi/IMYt8etIVzWNr/dZeU6s7bxPzpQ2kiKXjTcpLrG9jyALO8d6wHTkSibp
fe2XtKJO+HGgjc+4CpI5dRLpfm0Ns7rwYs/qBCdavG3jJzUh9FTVhv5NGY1qP2b4Lte3D7Zvu22v
EK21ipmj5weReG3w6UAQp4ZgY1bM55KMzwywqqpNgOJ0SbVkB4W7itRNT+uImZvvIXBZde41Wxfv
05NSAgsxyLi9F3Okp19Y2HVnU/xRY3vUTzJEZHb+drA3DkbV9KyDHKkpcyi/mJ5HLPGgnhifLu/4
F2Qo7cgR72ieCiqG38PkrCazShGAtMsM1Ld+kpXj9LcOz1AaXs66xmDMo5RN30JiuHNxTrZ16sA3
iUWtMiLIr2IK9komUTY5IAPBC+fgL/n5IN93xMq/5mW0HKAw+UwKkg6HKyMAd38pwEmLT4bnA0ML
UMVdAyJ1nPHZC0Dimlo11X5j/KoM4h9N1UUVZUp45nSn02PhgC1r5sEG788+rwJRaN9P52DuLG1q
UbsVHJX49yfyFZSImcTE8C4zauSk7iH8+MOiKBiIZzzya8IB1UIfJ3Vx3AKaF4OySZnoF8Y6dUPE
Ri14wQReBx5t0VjPo1ZgFkA5bbouKH4rD8I3oTgt/VgnhBpcyU0bJIVfANF4MdBP9w6uhpCTLsLt
/0alvlxzCMNEx/06HQ9F5XhGfpOupH9EhAZY4GXZ2k9QBLiXxDGLH6tCesZ6mZxGg3FMFQXhfFLI
q9mBeb3EKPUvFcPf2AjJw2OpWmPg29kxE6+d69ewmWPn5Qii7JruSpG9nnlIGKrtet89PHl4OJlK
LwUynK2wsHSgDCHFnSstnPH/NaObj3N04fMZ7R3hBrxgOQbfc0KUMjuu8sCL4mKTP1lqzdtfwQTz
MoMRZXc9+rcOw1CmBNo5RBCnz03oVyuCs9et6HyuJOWJengownFgvXkqyVPr0TeUr01Sw/RUGlY/
KRXQcXCAQkEipT7EBdag1hv5nA04DyJ5/5AqQxr1asx4T+zthX/Yog03riZ7a5MDyXaGA2kOnqa7
McT9MBxnMPkQPSSab3J3IVerGfw3MVmR1p7Cc8l2EZBh5b8NiFcH1v4LvbIinZjXmIDMG6d1Xh/n
yj2ihH3AMoWDxQYCxC+Ro3FoPDFFKPaGqk/9dNqZIYKPtuXPwTe6kEEVC2zasdB7Boj2c7IRr0A2
WwWess5zVWj8Qy9qSjja7zOPrgu1Qu5ZOSgGzyp0UgR4grrk4Z3tYQqpBngNEqlmxJZabbJ+Q59z
+Hbc73lJURjUYwK1jKk+zS44fYPXS+QWttOQGfy3yUPCB7ASPsy16LMY7iFyFOZQekIzWYgIfgGi
0eAfNPy4PRJBv6aJtejytMoB2QdZhyoa3a+x/gm7WYRJy/z2tMR1GN1Y4U4NaRL7wBx0Lz4HsB94
qSqGyCNtScWc0z/B9CJiffcKhemRFWgV5ZtFlBf3qq8Yg9/aA4ctzYID9QUMpjeguU9bfKqOPjhe
kW8DecaBV2RTk7VkSIHsHYiiDMBzf/8+i52homNGldUZq4mua8Qr0mZBvfKum62/LbRxAVjs57MT
XJOtcJRr2HMDZQMWye0gw+WPsupehsWT+Zsj7PjXlUyZlAc1hNJzMnmDqIlF96/KSGRcwGs/+OiU
rmlpNUF/8A+427peWTPWx29jAOIIhMYI+kJAlgqhi+CwfwcKyY+EpyVxIsy1KYh6mS7vzAYOBEq8
8PDDCR8UY5/YRwkMUCs3oOjJSK9DlBAi7i1Lf9XP62WBQL+reBjYOuJ4CdbzydfvTfFqDnsM6gO1
swP4CIpXZszy+GIF2TRvoezrTCRxZQb78NtqznhyJed0TU7/yNDLpTTSlRvuy/2qRMXERkNKe0Ei
j682HvHepmGasr41UIFmJLRIrWdftDYixDyxygHBNoO5x2XXTMj9uLtT0CxTSO2htLJuhelER6zR
TWIOK27EJZlc/EYzE7TuWdbkZOlp9nkw4KagEl+MZpC/wFVJP6732yq82aRIjrUbktpq3b7Ln922
iNsYZlSvIql90QUbhxs3HMU8rceDcPVIJ7C2vjwoTSNADoDtz5D/YTW1WY73qqC8chXTZMB5Kztj
75fq+os+bYuQ7ZszmBOhrzxO0YSNj1wUUSyN2gRULN2mG+mSoEfkqG8WAQDun+Yc5wdiLneUWrqD
XdiQ+80TG3BUIaM4yiopPATN0Uq4q+zi5jsYAfc+l6xTKdf4hG8J8BUJR786ipnC98HwMfJAEHLN
5UOitncRgk931N8UCqapdnQiFMIbqcKK5n8lUoPVGNPTn23kBcWAmdDkRzL3KL59p9RGns/S8i8/
T6D/IbO5XBy8vG59nByN/wTYlLgeDy25mHRAZUvY9q/BDoADFH2BVNJDD9luW7FGpddFYeOzmUDu
cu4hG49xMnvmbG3XdJqD2p0ZJhR4zkqKn+VGrmvxputeXstX7nsKkY4pNtAS38yfxhqUrgmOQRd9
Rb+zSPkiDkxF8iWceICPW9EeBcXagfgrfOfqzzX4qy3x9L4TFhsV7G9GFZIiNmqIvhREMYXiI+Uy
C7dC0LwNkAqqjCX28MswwxwgtI+AHFK8umYiHgCRjwPW2mkI4UtNCoWABv7Rr3oDGMIoxeoWLmF2
gXLNsoBfraMFX+A+9XhDAHVHFdV4xOuR1GhZyiDpmVo7eBCD6/rNJwgzp62QmPnVTdZiL5KLOcsd
tbUD11enkjGQ85bA1hM2KRD75RVG1i8hJ24IKV5HgCqKOO0Mca2QuFwdisGbEquee0UwMDejbPxn
W2V0Nc0Sr4Rnzk5ASod+X+MYgXKq2d+6NaA98WmGrdZt7ZoqeFyUiHa6z7NITbuURvAPToohgqpb
j846Ksh4oD2TG1ON2jsik/zob26nUPk99sJJlCuu8cULYa+vuQbp1KUZ0iIN0abkcmfRArZ26drN
owyRZmm4WFGYKOO41cGMfVV7pui7k2gw8fSeUEY9UM89w9gtUnKANJglRVvA2ykj0D3Juu+BZZea
a+SmJlGyNND5gOfFtE0eOaRILdp7EuJTAZgtIz23o6tBOWQwOZvWOofCsD0C9koPN3BjLL4Xvgjk
YPZREbLwYHe64It49FWPh3S+apDF0L7f59F0+bkZF0JmENGize3D0EKzQ4RCJPkU2cfMwOsKjtvb
ntqVRZO2aA3hsGjDSSR3BB0IrCeIsCl9CrVjYz5kvXSfThoI6MJdyFK00aY6hfUsAQ9aaQImjltC
+Wz0aNRf6ueocEL1ohIuQLj8WX5oR/WdrOm/78gSq9VJ9eTOuowrfLuS8uZjcgNK1qOZ8nkdTJlm
ua4LSBRobzifGLMEAXm4zqemg4gDqDs3FetJ1nJvG1voZm9GoJ8CJ9LmHpMV1L5QjG+USIw88p8B
lJV/knW/OMWDqKapji/hwKSbcWR2WLqgrpL2u97N93J70wl0Pd+h4w9/Zh6WiQvrWfr3jrpP0LOf
AJpn+qdV2Khso+tVD9IyiYL8UvNpE5zuh5ZIqBR4FtYM1sU4lhRWOdMBoNmJM7iwl/WbVSuS/oLH
DDiRZ+TaK5rseBKhP3LVdjENZXqbPOxR3FtYjrzHHAg1ddOrSYyW9B4eF799P7PEzLFc3GFBjF6X
m0pH0X/xhk/BhR0y9mg5zl0+pFO/FoL1XnzCWLrtx4P4/CSgZB3h1s/zS7eGws8o8DnBO9JyKtRz
SIabvYwvSi/EzHuz+y7iAFLmFGZZSorsuvfqZ8rZ1XWeAT4HFdP45vemK2Iv7FW2roLLe3WtK4x2
bQ9ZchunIxoflHBx/KzykeEGLuYcf9u53wCvkNV8hkaCMj4fJB8p534BCkGcXw1HlqDE0VFDKhqs
9RwhGxCAsQ/M8d9dhNUO9qYPDr6JcGUDfiOSWtaganXmO7+vAeVtiu4q1Yopat8Chr/6HQI1nLl/
Q60PYxfikrzA9WmUDPTlz4H+srf1sFjLyq2ZTBVPsYV9z0OjmAa8YsHE1cJUQIs/KZNv34yfKfRf
LckNCtLKdKlVZM6NFlaOJfgbj+/vOqzQSAcKz8UYgGP030vXjjK2scItesoa5tBjXgUggfYT7hfp
ZZU+VAuG9tR/8qg30MyqdCU4n5X5Vb9ZdT1SzHvXhxN++gUKZVq+sUyg6ETDJ3eyVyLVcnHtNWGW
Wb0QleQJu4TEukV9XYwaHcfGVSO5FpgwJpbqFXAp9NCs7P11EwuYAIMACatOonRIPtnADc5cF62y
bAruhjfD84i79I/JuwVLcIGLUSr2CSuFqwr9C+5D7SkEp3HlLd0SpftpOI5qE+/Mo4FuN4BfSJ7K
z7AylSH9brUE5AW0b/2TB/xX2ewEHW8FU+7oA8T7e1fiNqsXQKDiLgw14hhh68WgMsBJizr72h82
yFjLkRO5OE8xYTGw6ZeK5irxJhiAT4z8UJM0JcWZMTenX4gVucJPareZ+Bo9ju2Hgec9dluvfbAz
NMsQ7/HhOv+J/yKf/ssoQgWpf1yULKdlqRuXHsMK0Z67nT63jUx+0Xn+paecyqYoObbE3sXuIwu5
kZjPnuIlyD4jj+4stCAfhwEniX9blu0ZRJQgVIXcH9xtNSAt7UrKiDt5TFmgHJ8GnCwH1LHIqpC+
NHc0sH+bTsWp7GFMMYqi5/+1+k7JaRyEY8GhJvxFN6OkgjwQweVblnCaUdhDCv/lIAwlR34zxm6F
agPquSVDsXHFnxSc/kjrFvSWQ5ohUbJFzGodvD0vUxyyV5x9lktI3HoZug6GnrUE6DSB2uQw+icX
Hkl3AzNIVXY0IxSrTtSLG08FjbWMI70PkI3RHXKoCrF0yoDzwVvfzMJQPhaEnx5EoadvQ6FwnOt1
v8k7t9uObFHRb7+J9Nnsb1/VYfA7iXFd1ajWrlcE9bITYU/LZHj6KGCoftS87iFydbvEiqp4dJlC
9Z+Ah4aINFf1ctAPYoaA9HExbrNDs4Ofw/ispSf+UhJ531J028tJJ05BIiZm1UBpPWOa6gx+YJlc
6xJD+ujjXkkO9CVyocWbAbIIAUjeowIqatOvyQ/YDTCS0KOz9/d5X4oKt9itfJPjTSt++2BgJpe3
Hpiufj7VMPPIaoPYhc9usPVq9l1XlV6JXe8DRaIOxlR855i8M9mllv2ifGuftGFsitH8YunPZwUF
DPQSeCNtv3X1D419PNH/lIcTkCLXDKsRFyyu8ZAzBVmRd6nLC3iNNx5UfllPWWP/d/WdTNMDZ44y
l6ne6TmaTHi3tGSAgAdY5Ku/I2T4MlEeJ0UWIBtIdj3YbiEq2Ny6EpojWRkotefPMit2GfvjXK//
+yNb+oTVmtddIHd/IRZSksw19tyMApmORlr3uDENrlKkptOg9byU9ZTzu93lX0ipLbqkt25Wvd3L
s+PWhiqOgoF+a4GEbIFpE7ks+0JUzlyxGc6C+a3e42oxilcCvolejSR4iOig/d5UDwsXw3wqijRz
kon7/ZD2gj3CNol9FE5ZG/rAfqGO66V736TB6GuNa6I8SbWlWfLB1kmhVxeJxlxR9zIr4Fl2w++V
XyK56K4bF1yvb124JaXOFemJ8uxCwA6UfYWzqSZEfRbotdpcpEUO7bUYijO6XtQDTujto8ggtcH0
NjP01gLK3WbCKvt/omD110nRI7ThK61ti7NsiS1oVZMQXNwjPM2AqcrXCz9PqkP1Sj+ZqWXVykSX
SKwsRQ0IC1RdhMSDRCsU/1Hn/AekMMTrIf1aHX1DN31j0NTLvGPV9KWNaZCWbyy//Ad1qF/IBZ3r
bGUQjatrzrOifbsxqBv+brqw+a5jUY8RNyLv6nywZB5Ua82O0P374T1LdYV24hpF0pcSuBfAiNM9
TuuZ2ZcJNvIy+9yLiwv6gGf45Pc7eOBlOn1v2OkzcRohze0uF/I+vKTp7Vj9wIL+ZTMz46fEGa24
0vz8p8ceK00670hrctuorLMIuI1Wo9hzK9J10bQ8Foi1kyTm+QnE4hMDu39P2GRTH/haHfFy9OhA
BNNK2qL1GpZEDXdH7kIzE3OfMRsiJaykmAfQN7ChwbfMb57SI0MR1B2PzkRA8L7xkZRYLHTg6wM6
FN0RXMb9fdZWHmTDAHoyU4O9MoZI0kpmMzVs5puSbkpcYCVwsqbpRo+X0Dr7+JXWUiOiDZr1pB0J
q2J5gfE3YtvovFXNhd8aBpmA/jgc3g92Z2CzbozgH88tgYdMo/5AB2YM+NJTZHZ78wmh5aLfjWRg
rKiGq9HZbkKO56a8wgmvRe/+SxPpfUvVJmEJ4PGooAieRPIfpcmPno2KXCdYFiRYWL4/o/OwFOvA
sEOX2wzYAKkeDa0XoyY89RcoCndpL9gIOkpUhmOPodivNZ/7eh4DKPaknmKne3XRcjfGCV65mLIb
03JqEP/jiAk1qLIQOt+vmqWS/U4spcR9rk3Y0bEYSE1vqFmcyR42w0MzqyhZhaHLLYRUdJsMZHmM
CdRwtkz6sYHLcfr6aA/BBtkputgdx5PHaREekCQfrA2GkMrfQl/DrLgqGvQz0PZjS9dY8k+9Ao8G
9RGcq/mF30ljDKh3orp8ZO+GW5f3OgptC5tM35vSg35TrYrJZEX6l8Np/VihrV2/8eF++hUonUdS
fwzwfSbz/pK+C3Zqrf0ogceowEGeUZKOkJzhp5sh/YbKs13sQihKGhUpMjpTCJJVpweoDjXZGtuu
MRGW1EHIfpw6WTcaY4CAiFdAc6eMy/QwIjLS+0XOdQMPph1bW5nUpLOFKZNnFvQzFJIvpl4rBU5a
hepMqe9FI8UVkoDTmplFA6ltkzmYpNx79XUZPfYg1ah9bmk4vpELmsaj/g07Dj9s3uumfvk/wbqg
Ndcf4M80v/A/9B/hyPhZui4/sZ3CFLG56czhjr2MiYa82XEpqAVjjx7XPmpVY7xuJ4ZGy5XQlof2
/7lp+vZWaShQ2TDc8x/XL7MoMldzctffxAr6N+X9FI9i84w5j0bwG9XOhUORTqCUfLHRgIxaWC8c
9k0HBCWcxaNCqvcJZyEI7FxXdv2LTqy2gfFSS7uPJb+vMKTmyP9lh1HjrRI3v/HAtUoEotLwX+7s
M8yaxzTVxe/01dzwXcAabm6lW3ECe42CtNSDUiUNLk8TEPRMZOscckK+zWIQLJhLDfJNxGHbx59y
j9/KiWpGe7Ehf98bMvJgRwdRqAldArK0Vy3o0h4dtwP7ypwrsUO4UMUSnqMyJoHm/peDQcu9EkGB
PR6z2qMzqbsDyCcS8B7lgR00Tt+2gbdfZtYw3Sz0UaRgn1gxmC8jvs9Lobijy8efO6t7SgiPhDIJ
cxwu0XAgTyB5yfnEyq1iFJPvpM6Meelzw4E8tRBgjlNQ1mNmJkZ2jl9cr1A6u5eMzFcVhxTaCGlq
04sHGg4frt5ADfDz/O+QYfwS7lD8o3Jf8tMo8Ek9xnKEBCpAu09het3xS4TuWIhkvfrzY9q3BSR6
bqOUSTlHl0k+TLo6hKMeJHZh9Xd5a0GxOhkPyaD6VLlsHsxnO1ga5YEdJjf0jrglxRITxWCvdcTV
5LVomI9XdX+h+GaKuG3n8Rqeqv802nLZ1qnYfYIDdbFullaogjEwpb6N5b1X2fygoyvXEHAMVC5C
P84gJ78KEoatfuPfA1AkRi4yZ7JW7tknhm6nHfdeHHifW/dKiw/c0QMXlS4XLfZxbVRcvX2au+5l
UTdOEgFXQhHFLvJ/tLE4+z1UMzanEOhVOhEn1pA+YThHSFr9KhJFy61BWW8yprMHhLbPp/EiZaJy
FKG2sEU07vDX0SFM7AoI/RLlzj0S0+FgW6nMcmwRGUqp7F96HSrxtj8kLC8iPX5l8doHUTLnG9F9
INeDRLp1zJgI/pTVTVuBWe1O0QYIaDfD4S2fyOB5vSS8zeBgObuhznZhA07Ow/fqP7e9vnkkKYVT
O5xs3q+D6BNTP18Hwl0+UaAn/sestQbfJYvnShsVX02NjJedsnCOKxeVXJYW3LIj4G7aK7Bsf2Co
+X5zg9DlnDWe/KksNZ3vPTAV3CVS4ovHwEX59t4D0DqHSu9DDaHEE5ZdTEDmJOv2fZAhbXzlvnWY
XbK7m3+Z0rtlTud3+p6T8YhDgtQQf2tvhLU3NG99D18bbt/RKqW6cf1peD9NLGph7gkWDER/6nU3
Tj67LxxhA9s+B7KwE/uRbcNxsRsIr57K21TnnsoGpA3xiJpz7XpVu7qn9hm8Iel8/xL3gg+PkAtT
YbJoIo/IRk2WvSqUGQrcSMku6yUw9+jf8NZ+QoiihNjUjEjPMR65XsjH59Q5KWRRl6ttvaALKEeM
l3gl3S/lmVfYvmLS5ziAvpijxfd75t+x6MIbcFqr9V9pruUfmmUKMD8EWgJe6EGRDRDqsgngRjnV
9SHsqJaJqI9lkpYxV7z54zZ06aKhTSM4ckAYomyw0jERa8YpORwV16qAG/kYVuND5/Lwo1I/hDum
QNN6iIRBN6PfiqQhv8ZA8FYSEmFYq+x3jg2ZzcGoNOlCyJZb30w6jWixqCTVPpUh2qpLm9zTJ3NS
2jG08R5T8pgwLTqfv2HDz3L/ipyPvGwmZIgbqJQSfBq+rc7s8bVhHummq+KJzu7mp+ByP4T8xhAh
taxV8o+IS1Wr6mYnJq5vhMXixqBKVXYN6L3TlP/6sBEPdFboli7oYy8s2zumJoBgPCjYiRIDC88Z
GKnvtwgVPkrg0rwjSI6JOt71/G2EGYk/3OUs+2eVcB/HSnczCavduP+7schJW2G4nRMLys10X4gj
qLKv5ARWbEGYwZ/zJXV3GjSw7fnBrPz8smKiwokp/fJcHL7WIrRd33zPI7XOG9boyutnzTUethFs
RgMf+yC6E8MPYk2Lu7CGXODhVQ8rgbvrqdzCaxvjX+kj+T4IkGePYHT3lf73oMfJNcE9KuYOWyhB
BUSoyQhZbbOdkP2YdsfywjD1L0YLm0rtM/sNlR8RwWAFHMvA7+ENbyB6BzdkPCmunfzzktGMG/T9
vmPUzBm6ZnL3lmKxW+U9jfs1N2QSFiQQSPMy+I7lNwwtkh3HcZv81uzvnUMvdyymDg4s0HQk1aPB
fAYtdmjJdFoDgR2u441rgBf5ui6PtnpKNaqqGGDLx3LP8BN2dcI91PWwE9VpvPU7JpHyUcRH0+Fu
kKGVxJ3fGimIwJGT4H/EilVUAronp5U+REAZbvBzbJsgYDxpZ/Rklsk9fkO9g66Bf3csJ+clQ+5H
w5r1VZtZdh6nJVEzksp/Z4EU9bqiLn8Xi4lmNMf4+EaI88B1r2sdL4zCs5KqQJBIrG8g0aWIsHoP
GZfkXxZzebKBgqjIaog2/+YN0ka6/uB6xsnxr+A3vHmTThKXu2Ln6YOeqVx8JBBNEtPXPWLIIwbp
9Tr2e9MltJdJgqWxnuYAuJZiFD3aG17zms08RqXDKcTEhZbVGdF3tvIdqw/HkAa0TVLltDzd2sHI
EfJQiZX64AavwEhCDo0+42jni8j2gZrgGKiz/Qix/yrwoASvmFv/RszDmLMWiV7yo1nQyaaLDfhM
rIBY9doKWzj5G+AakDruSEhkDAOjalhyHuWlRivZVgU4BXhz9rHxHmsjWQ2JzKwbfRPoIlJDD/54
nCn9cazD1LdwQYSs8mCwWmpFGIYMANME7GNwkaqEzEEt8EdN2Hu45Bdax4yRRPtECNsd3FDJ8kh1
oKneEmsIIICMCBuIpLTOuSDu4x6MLW5eSs9UZI3xoqO0hF50m1YEVK5ya0l8OzXbz1vg6CNGED1R
JxDVqbFh3iRToV/YSY2Z4HLTtjTOnDLrmqix+Em/NE6SAPh6bp+6hkXzjiE/O4Q5kOLh7joYqXna
1hzjBENLrPdkFdEzJjOCCUX1kERc1LDSNenR26A4LCG4Y/mrVwS+wxt4EfrXtYemi94SBA+oDzlx
e0MBWtCfBMgrGM0/gX6PkHUfa/TrtNzQoXCAZ3tpa9jkAj5hx5XNyatJzfJYCpxPEnUjb4Yylj2U
n3Fp9jO3iireYhrL/y2LaRyw1dB4IbYuXoiYw0Y0djfE7Ax8Ka1ogZeMQQkk+jKbpiBS1ZSF7yQ2
YdvPJ2StIpoQALu35dD80BPrHLTndi9BampYhyHbrthdiEHf9fUZw32feIaaWqIwgVNC94I5MJLi
CCSUtPcYdy8vvoeD4ShsoTGIA79et2xnIZsWHLQNuxKjiHJhEknjLe8wc/f8+Sq7CV0wQ1igRPKc
nKFW8VtQGKBrytubfIMujkTBm5zbc/kAGqZEqoml8O7no8UX6L8WHrQLK7wMRyRBqBe+JsQsQW72
c4bD8CZyy9PgaOZMRTw27HU/dfEGD4NXcPPlJ6dvxRrQj7ydydTmnYnwah15KsSMeD2nR2xZYbyh
N+ttZnRob/QIwifbiPTzAYH/8QJ4+9zQC633rXcfRJ8uJQBZdXFTpgmUeHao1E1MyBXntY1Qf+4y
U9DYpYqgQO7cxhiVwwCIrgzL6fmodmmE6wWTWTkbCSBzv09+pjSe13CvpmV1rsK7YoJiCo7XxCFw
Sb15tANZqdoNu6Jm1R2/3ZRXWwOLfE/kgwat6vgMB00F0Agj3aiH63P/5yQxbbITEUjnTpaRKtu4
2XKZQUvQb+BA5wj3teyYD++5oeFYAqO0kKvO8cG7sC6uYQLRNOP/Ie3xWMD6A2Hzb/YeFjCLrpX5
2I73swcY1NjnE4nA72HIuw/fxakKbxqwz9dle/As0NexnEUQGxAbBCgso9xAdE7ESMY8JEtpoI8L
jDFfH400bHR+seQDeK9ngEl5ywANoeX3Rmh1Ov6NcQRPznRRuL4v2mnjlzsSWUr6iRyMi9edBLa9
gdhGQoUPRm6jvCBQaoOD+v3+5Jm9PvpvwX9RAKsoNP+70zNGDAjGSwGr3q24jilYvMJVDgz8+DF3
kfWGdZVjx1FxncGA4/tcKvmu8XC5VvoboFxsjA57VqfIENLuX6Q8PsSIiLK0HULC7tFCfwItLsaG
EgSyI9fc32QpJTBb5s9Xnnl4ws0akfWBtyxNQhaXSYNjQeySeVZEpQS0RJ1CcOWnsQzGpQE5QH6L
8VliiQ6U4b9pCM/HbK/jT4Jb6AFfGJzDZFizCTFV++xRF/oB7DmkoRlbjDIyeFaHLKY2Z8YCny4c
3gZ3qm8PcEjeGIGcQkLWJu3lOsriQYqqwtlTZUB8cmR2AK1PvE+Zzj+OxLBh4FN2DzxE7v5qCDC4
T0tCWQbdnrluhJmVaZr0/8PA7NjMK1GUanb383Kl2PKX4XecG+jjn4nO+LzlJzTQKbk6W3RaPGus
k4nBjcxqpEQVV07qUZX1XNECauBhLVRSJm+TNoKD2va7Lv92gn0xhJ3TBVbh6USF9jkqHM7YOx6d
wsrXk5nQE/gc924cIiBhQCwhZfqI4tLln28+Uw21W4yeu+T5edBFDde7roPmWUaJHTRCzltZodmx
Vq45NQOs9MlGNQ/6j8a5S6BJRqDRfY2znz0xo3xyxj90L5jZqei9+QGjl8ME22nOzPqwvfbPUy6U
11tCPcfx3O4IArhFC7MGzVaEbUNmLsD17ItQLBKFRTJgLQtOy+nrTHBTn9Pbnb4vogTmJGz32GqM
i52EWuJnoPfDC/MCf0VQL8eWkabrnl/CjWISizTc9l9ZzIYa+56P2eQRBdaqcm4a32FiZiSpK6w/
+NtSZFQyp7ES8XA9A4mSq7kplrwaoD8Wof5vJlDgI6HiRMEFl9FBJiqg8yXhIWra8tOAXKHVjGnL
J6J2lZavW4qYh6tKWufiS7/REoZK1Vmkgztk1vNrTEgyY7R5G3RivTP/6AtZ6PKXjhhtLuUK0Ymc
yBaPM+1BIqGvND4aJ0L1TBeMYtZFhuwmzgUEUpNMHNlvsDgtE+0L+H6ojoKu8EgVK3k4zPI1qQJq
Znn7SLXbn3LWY+WFd1BXboTXQozec0y5Qt0FKSLVx+ThSEjRXRBqAcuBAXet2vZHQCNJmaZ924oS
lFC+WPbgRGT2wAT/w9M0eqqI7lNh69jAicBxReFMT43jSGADcp2HVI9nslCtIMasd1vqakD8sqO6
Hthb8bjZLGPvDfEfOrO+VcVD0OwbCEAkMfGYXUUyJfMo5OHyfDkQHObI+f6mgfT+E07mGh1wHWC5
fkqvD52WBgCbbROQ+BtZ4/rpfAWvesnvAbrKywk+FezlJdVY8hRXrSKUyT2fniqGC3dOCBUV+1Sb
NBlcu5kY2Dt4HAcwmc6x/Xa92A6O4ZaiZbold1eDdSUmxTkeNslULtFphDlYp449tm22I10pCIhQ
OLvshSNDSDQWv+s7EfYjO24Q+tkEd0xVqNtJzQIDdqCrQyzocxCbCbhTZBE20CZqpealhukscRZ0
lFns1h6/aHq6W1wVYVWYj3FguPHXhln4pGEdY+B5vHzoGfgev4qF8r8nqXiC6rha4Lfbglzf7QdB
WZ4ECUg3VeuEmg2IdPEmuXjqhE84HB4HxpGtxGQgInUI1B3YlVgcrYjvKNkwFPvdvsRnECJ1gGAY
knPVej/9cIZ11JmXweGLk55QlvjxMxrgDOm92gh99xTEuIxUbdWa9jkPNuNV4nmUW/wTpcsfjeGr
R0003oz/dbDeMkA5yMsicvZxy5X49S81UATO9OzcZiWePaDkR6rqAGKuJHmpzMPlYeW2MmVTe+3x
vHficYSPMYfiVoQ9xYtJS00let1M6mdlj3LDsCL9yhgi0Pk5iaUmt1BaSPmY6RN4/g+W8p9ic8hL
yJOrYMwDra36rUy0/knXFjZNNYelQC4YcGP+Kz+geybJ6j1XP+YgiA+Vtv7YCC8sj4UIdaqPlAq9
c3VRfDBwt2f3/C5XrUoI9DX2b10DbiHUwnyizNDPLrLUzudDV3NhELdbxq/FiCuEjL7A5GczTV+i
v/UoCg1tdQGTgcW09+PcTnG52hT5VoGBQB3vryOZwd3RZOHDQ7m5CsAhmhbrOb4fJOpyS2PTqxl3
fnMEKiD1mdTL0IZi+39ppaFmGsDoPWm4Hgwn6GXghNvnVG4W6635bOYeMJBunt5jY4cdPrCXzVCU
edgkUe2UMzHX5egCU2lE2dDq37K3B7jjGHzj/BUZEoX60SZju4aKkgtRVH19cCOKDqXLcPzkhVLs
jxD8enWsz8+1uacGqUkiihVWGg8p002mhyZkp0xhUD1yXIstWzPqYCOtgi4yrKWsKSe5ZBskQvjV
OiUMm3Q7Jrr2a8qg3vVUSBlOYJk7TiJJwHbvOYE7sMM/ZIBzmPQWYfwIBoyMXRJhsr+j1sAtDwLl
T7Nsidn8CN+ReZtfvShhiN9/RPworFNn/CMS24EwW1sg1BJzbB1clmeZKHixMfqzu17qemIG6n7U
uq/EqYCQL60dO9NHtnNCoWSTdSjw+SFCY2WTw1BYReSgmgN6TC4MxO9euA3e+yaO8lmTUFQljrcB
9tPwQdS/h/SdaSsgZlIwb4qTayMxfBOMfNhiLXiFlWBa/807jQbLHleMOMwh54yDPy2DzscXZD/V
payo8H8itgx6GwUtm4qlKFw3ZxAm9VtvbfAo5ztysYGpjkKYYEWztHW90nbMW4txUsPnmbc5nttM
lABJ87QBW+CDe3bw12XQsJMy0KBP+CO4ov+JC41yGw0XHuo2lqZ0TtQhnDO3TmNNIT9gknUM/8Ux
JI7iWGaqypEpgPFShq+BA8iBy9QnIcKBwCyZ6H3Dks0bP74r6npwWpTxG+xNyvYVIcZoZhibjAZB
0sZM/XTIcfpIdFeUNeyHZ5AlMQl7AYs0MICLGyyvpwiK4b8jri1Ts+iMkZAu/UqJViSYaflisdXk
ZmQiJ4f0nMuHIM+FCpZqM4zDuADVApAA3/NimayMpmCWlTvDgsQTv8BhhQM+Aq7h3s9opZDmzTum
fkvnG3e+G1Nmd2pObchmyJ43ZVT+9q1G3gOENYZGdbcN31jIvMIJmkFbEaHxlRUYxbBy3Vuo9UxO
pp/3pA2n30+FqjYzujO4xb4TzRL0yRrOcO3uK1gtrh4ZuZDqTViUbzL7Ki0ZdUVv2vrDv15Ktjhz
khlqqwpA0LgJcYiFF69JTJFH6Up9fxyX2bFooYu47gPuDd2ehY19d8uW5XzvPXx4oAve3WDGUQo2
SNm62hqH6qeNGu41quism/U4pYtrZh2KWSbd/WwBjn3rrGqxW1lHEUoyxgoOUL6E1BdNIyEHV2oR
6eSdzysCybMBu0JWE/FyG3dZmw8ZFxYTeIMtMftx5L4dcuusKahyT9yf96i+E9CFazO2IS1WFY8T
UiiX/pJ2IZDsUZtOSIbxDcbcO/ix6w4Vvvkh2HDNVE22DcfOodnmlH7A0NQ++2hXthELP80lhXdO
vWobUAuDBcYlGEFqJ4Mfr5wbEXZhWaSPOhrJqzj4ZjX2vrOR5LUPrR5SomGIuUXJH1hl1pqWtvB9
XuqsascKeSIElE3Z5em4BkP+7IoOfxo3vUQN/6LA7YV3YnGrBjC7pidI3CujWZ6qlU5rqFGCA+Re
+JpJHWyOihxVxNEBPs3P2ltLh50Vsm3WjtnJDZe+yYUOnFWNUj0tbmtExY6TEuVFV9Pqa4+1X9nL
MoU0uW7n5CFf1C4TeoVYdK7WRiJ7IeOk2QFhJwiXyjFKY4zVVHgOUROEsWbCggcyWSKDsAFfLgkL
B675FlpM1EFzuRDTACkWRfqVSSnTqHWszI+kr3zDqO6jQB5XxG26KVIuZ7ZeMMTsytpAfCQ1DT9t
dkhQJOzpovaAhQPHMOVJ2KiX6lCWzsYABwCHmFsxul5z0t6UtOr2BW8oa79qTu8ffgHdNr0YqUny
iM7j54ht+rQdzU3CI6hSbflxDsXTYmxH732ZIr7ZG7m1ycvSoBGskjIsQpBh1+x6/fdJqDw6C2rB
wCezWJwVqdJfO/HDOVVXbR9utwgZ1WAwHDTLZkvLpv+5RAUR6Ep90K9aFmHut/7zLu/anM09RKXa
eOajcPSxeL79tuIE1QLJEWihFvxjsRf7QgWt9MfojOX4rAPsVZESUqcov08HtiNYWqratN+9cbLx
ZyaPq78QPf/tWq2YoQ9J5Jbd+UkYZ+69EKsZwxHutx8Gb7FRsXnO+pU3UuE6WNvoLfQoMrSRv+xE
SQmEqLuiw3AkMMWuGkQ+8JTcBDZykt6KsAXtpdwtInQqGbbMYAIvcXyCV/BLCRVlc9TZ3Hczr5Av
wWavYSRgaDoAIEAn64Pb+LmXS3rpsGIhDEkV1XHtqkbFb++qx7YIB3x6eylVBOo/9nSwGfH8Y9zH
ms9PawHXQ0vYIAttTSsV/WBAQMhaBAtDWyuQD7yGB3yILRsx3kQ7ym9XbhTbaQ5d105jrpLQvIAb
DFt3yeQGWbHQy8FBcC7f1NGgXjX9VTDzFdi/YnpSeoili87TOLq0KTFAIo7s6tRaT26iQMEGCfEk
OCCpy0xVkwrI2rgHGT6ZGr5tEC2Fj2nYIS1yce6R0Zrn0B+gXhpgi/d0z2hetFrmlhBiEhw7tEAx
udmCRbUY368cW2+N9qZaE23I3EzOYjMMr2ukJRX08OerIwOx419Lf7SIG0R5MhlpzspIIVblq6wm
W/Lj1UMTXV5kGwvWj3UzxxritS6GisZQzuAkukz+iShV6B4PBgcjlht8G92kxaFxvRGRPswLXcp5
Ch1lDWdHrYFGwsCmWnLF8W268u0Xl1jLewtCSQ+bCRFSmv3jxwDVXxhrmWxD5M+V/RzKXs7hb/Y9
6U7qiKCtzdrWJL6g/YEZrHyw/YOALDhcC74+qCm9+FnJHNX/zpkT+/JscvAiah3qZHfBMLj2zhCo
lRYRjSyb5Wmp6XxBbG7OsR6w12fqdBp/hZi5AnIGCpjnLw+04dRzZsjr0XC67x/f7wAWqtQE1xMB
kiVu1WTPLq+AvN4ecWzQ/h+TwYlXmHKhwyiYJtR8gytwjnVMCa1Mhqyz8f6tWDmXGIcRZ0umZMU8
c9uGzCWEmoAobMxM/+sFBB05mSGypldMphEhfHPOHiAHV84bnBKwIYz5DvF9ifmGE4NgqoC2Pn1S
ad2fyaIy/YdNbjya2/M2dGnPpq2pSccX/kz1b9YZohNBcYcTCLJ1LKxZ6B6RiDScZSj8U7liD4Qt
XiDg+8wuLgmMeEtSNwjP2pOVQP0KWbWXPCtqtHsYDGg/xFolUCUCAOnpH77ro0YumVnYbPxvlk9Z
3JoQixFvvBjAXnEXMX9aMdtsUJQGaIiOcYGMtrKCiRNkrWmuOFzFVuprAbBC2KVDjjYgZx75WiHl
S50XPeAl98UKLebmtm1ojSC4kVX7WyTzNTr2Oj6JshhWcvX0zgdYivP9eB5eKNOytHkBxTiuH6Vb
pIIfb9qnRmDhw66N+FDLK/Ypv4uoAJGfMKc0g6aIdBi61YXQjptVNRqTWreDQFpSoEVdizfs92SS
AgovJQPemlmzgHOXnFMO0CK06V8Z29HtyBiBimosrhH4Epra9ZygqDyQI072MFJO7/y9iI4A8lwi
ssZ86r8PYgQTNBye1UJ0LT5X30XP3kOguiMGO3DtHqfuIYAvRB+COtfMNNDOx6WgA4pa2KjFXO8f
eyxVUlhC+CBZdHID2PyjwZ4OFpWFxkZ4f2xKFNQPRogmqSqMpkHmhqvYkT9Vlw4SxIL5oxfq08s1
WF6SauQlDcjD9M9QccLDum0neiGxr9lh4/k8Bkx4Upnnv5Zm6rglhGYNHDKiE219N/QN4TIXJm0Y
qifVpnP9P/Lz2CAkxRLAHojyisfhlcI7N4xP31hvFGQ5TupqXG5fA6+tfV2/FhgP0Svtzlmp2Mal
vmt2+5eS8lcDYM2IitVCnaQhvXcKyi00xiQgS/EUHbaKfMYqxOtm771dijJyAHQJiPv2ANIPcPc4
BRHPbSIBJF9sUBK/EbQJJNXtLCM2v1Qmk9PFkmYhz0GRPNwyVWTgqBXPB6vNUUWM0zuJpJrWVPuw
CL+AxQW3AJTLTtSw0TR9qfvUq9I9UXmm9w5ACEvtpu5+dospHy8c/xGc+gOtukS/QrVO4mmUxy0N
CuDNRmzHLmAbBd7CFKgWktSQ2tvBVVd1fnSAl8PBhXHIMP8i3FWlw5vyR/GeXrdZtvKLQP+WUBLr
CmvNOcfjpKeU11kpoe0a7un5T6yxsDyqbG1aDpoAu/fUdauJPUrJs69f4+eJELb1WE1mdlyY6W1t
HBeDRZsUosM5QMHv8hUVXhcfhABtW94HZcwSuPKTpElsiD2lZNERh3tYTQv8wKEOCXloxgfNSFBi
xIuj6N/4ZDffMYbvJ7w3oV0pts0Ro3yJub5XCO0pq+V1ySpxStAZKUWCg28kxSFP8baDx4FFYwMI
d/qDVDc9dCC8bLtbw0AJ3DeHxuGRm0NqftrGqTEpyTyWIlI3PK3l0RARegUEa2ePjw5ydDJ+x47m
w0T6UpJyQ82W94xLK2AIwlmgW9cKHjiqDGEWpPkU83O7nGoqNf+NhDSgvcXE5cijm2kzpPE0H4Xn
l0vQLZswi0YM46DTAbpWRNtqgECCiXNhDhrMBXhf+YFemQRYr2C3Q2d2afWzzZ2iasjQu1q48Z0M
pKHak5yaw8+CnsLRo3p99usxoYBYRTqIRtkrvIHZQ0AxNs6bDYnW4M1HX1cm2bpw6eqZp1IOn1aB
HfjRonoarpbRdQfBa0+HhM+pLZ5q66+oEg3kdYwDnbthT+j3MgAw0CFHPWohzV+zBUySjLPi73ZU
Amm2QIEtV/GuJjFF8aSFbwolkyzWHa4OEV/hiJNmuXRuV/8nnm4lW3+mn24EqaOjRm1VG/Y8y+33
lBLJoJNaQLjk7MBqVsMc1jWxDlRNh1XyTZFU1gBMZHTmxWsksiInp0WzRgvJGansH3jbZibwGg8b
6AtSJTKwE13uFdR1gSyDpKu/jPXVwfCU7D7v1fDmeo2a/Bm4cDUC842JT4mwRAkhFtdJ4P1F027O
9EJcnVEDO1oRAqS797yTO5HV0IvsIDW0W8yToQllReHh7+n7+IQ1CKnTHOX7qa0qiOw1mp22Sds5
eDDBbTc9uNp3BZNjm//07I1N1C5LyC4HWUf/N2dgCpeKoKam3FBPzhElxkXd17hlA3cIaRwDJbTT
K10K9FquLCuY3L/PtRgfZCjd927pQBpZ8qMhU/T27E0PbpwOo0YueN0t2Rrkf+/D7iV2yp4iKSfZ
mvau3g1LOcx7aI/fqRUNlPvL+lnVACuLl6FxmW2yFgdzaPJgmYWn7meqT8v4RA7AlIeO0NmSmfwL
jy7jWWSFxUcCCPsXD78ixpN91MG/iysndMbbD/Oim8I9o6x64D5eVuc0QouPeonm2gfbs1cFf+6N
qfFt/zg4/R3xP89WulLWWN+rhUX3kmBhHW4DneIQENhPg9t92E4dqC3RpOF1U6x7GEI+8lOOMEkl
l6Yuw6zMMDcsY41KXpvy5Zk2yrk7zerd+lAYfdg6lkjjavztB31EQYis8eaCd0tbFMGGVEKnnyxY
zPHq7F/1TGnag2a6orjznhqVyozWbSmAKG1SFE5+HiIk1DUlxJgVK1xF+RUzFPjP+9Ac79GtJstr
0Fw/SPkvP23Ml+oN6F8ohhD6rfnkJ/CE68uaWpt8UI/nNhjRLFzSKTv4gwpazPQZNsz1Grp1kExL
39LkuHElo7Dq4jEVdR48NwRZQFqm/dB3nUiByTiqJXTjGkiDv1HMmOTjTDxtPw9fToGST36ay/Md
o2SL075htdJEEdYbzQk18d5W7vJZzlQ+H8sA0swVYnfG9zgdaxk6S3sZsqNjMk0BJcEaUNRe53hA
fYxMJj/1t+0L8L9C1orUx5/VLy99JlNbV/92Qscf3YhGE3xN7oFZHjImeg2X9KTQJADxmky053Tr
HXxjUglHj0tXpnewDYtBvkS48sC63MvqJfMR6+QK21aoOFM5LuJuHcvtYmDcIHczvIISJlXyDXAP
0MF6VLkBwIF76SSYdo1rQpLDR5auVPtrJk2M03rgTJ9WGNP+JaT6mOBGvLDQH+9D4EkhdLOsBRWw
TSeMWqJvm0bpsJXnouAaGqtJ9QO3p3+WOqUEWOL/coIcFBGboSjhxoCxrthLIZta2c5dOfHA6ANu
EvY1ianmNTyxZ4HmBivhHSLWr5cKO9wtX5ZIe8V0gUevaj/wcQ8tR/ITcIdfmECXEUTH/Fvv9++f
ziw+FaRO7rDgT5rV55+RbOEZaeMDibkIOkkELYziRyT1gpVY+XR3aLnFCdFpSTjzjdOZzeTQ/SYD
neZLuvpXIU/wOrRHK5GM/iBs9OCMr7VIZv1mcKH604G2oBdsyco4mfXCppyZihxUH/aDbD0bbqpF
dEtog1t+5D8W3JXUqYTcV/KMYv6tz3NU9Vu9ScgEeAX81IT+JqLfg25STdCglQzzv8+No7nNrTTI
JrN32jFcGgrKfnTaCYy/ITkQweAanA+NLEjzjaUv1t+RuRoudwQaJUGVV/2eBcoTYRcyo5GRLXQl
DE2rtOVdbtrgPsssbDrVZYtQxaFp7XLbLPGd37HhCbAPFA4U+pD5omgxDkfRe+a7Es+7zlE5ZX/T
ZxiTVJmKsl0aMr3Vn6LkwX9weKLKI+W1rtLcsF/UE63oKPLVaUw0lFYjZwbwtKG2xsHdJjxyLqUX
ZNqDNRu/HfpFKOhQm9wYgW7G9qRTtxmxI3OpV3e/Gb3bgUkyQ/sxdfzVe9fD2wSNQtYwUSUcws1V
oqRYA3AD/jDuuXJ+PXlmFPDfzvYLtgKdvXkvDn6tbdyYE7j9tAz/da9Z7l3QfGBJ7CnDYtsv6CNa
PbxSXzXUWanG/JHiT+Jfkdp4P503ukp5Xoz6XC6POfMnapc9giHzdEEsQCQixm+5VQE230Cxfx53
7mymnZPlZmTcb8P285aU7BCVNhAKAXbvHoPZNys3aJhrwYiRtYRRuEXiybII11rpAm5tf+3uVRPb
kFQ18KAbqcOOR3VIXzDvKi8W6LRMve7SHaJMhlO4OiTy1Z/VzhydZEXpyL9IjGEbrhsshhVeGVAi
7z2R2gwecnlFX89f2sJpsULWrHM+NFH0d6hm0nyT8GWzB3zZpVSojA0j8spwFrFemPGZVIGaNNMV
MWWGgn93MwBrdkvyMtJqqveSBxaIvBklNegYDuOQpmd87FZh2pXbJRKSWM6z9i9Qu2VRVU15sSFT
MRA5/MhksQN8rXDLU1a4ryeZU1plyphsydiwowYb8HaUehjbBkWOHFo4HWl2MFdhaSRt9odOjF5f
c8Lu7qyUHNBG7mJ9E3qH2+REMvVUS5bZ5B2FHN+TQ0VXgn4oYlSitWdgEoFWdVPsT9b0OdIqAtb9
z/eluxW2g4beZvvbqMB+ORLxtlrWpAt5OmN9ds+4zMtm+PFpqcZAjFNf09SkR3SPu2dVyA8HDArs
DMcwd1HagGNo8XnlMdD2tlFzytTnyS/DRTV23Xryo84L5GDLRO/iBOmKkSslzkn72OLuVZP0fNTM
2Io3rf536VmSG2J4bL+ldFD0uf4p+2byNZp6mCDgL8Tk9Zn+V8XWx/iH8DmWXLKyIjW9Ve1v5k2p
zKX2oQOCuCQpGyvw2uAWm2BFxZ3GE0c4V72SaWpMEBfzmP1diOEW+NE2+DOavBIxi8azCmPC8GF+
wJva8Io/VgiO+Yut+ShP7+6HzeQRTuOHcndIFgMwoZWXiy2d8y7yycekbdS17PHcEWEncM2lZjz0
bU0Cvku+pLYF0wIYZyAgc5VGhKdGHjOBso/TOCUoW1t0frU7sAimQNA5sTzx1ChD7SDErBDztgkM
6kquafjfyMM6i74vS07w+sEASqHOQxP2v4rHiQWuCU0LyeIpW2zfyTNlL+1XxI2Iei4QlQJHqUYc
sGy2YpmP+72/rFV1WXGs4cwmsPrruBpMDYiR/u7uFeMLd4lVGhrBkJUKej6F9Ay83LlFkjlzqiKo
FSiCnRJDVFTKTy6JSL9abATxPYkw48dfNZ3dCI4J11EdAOagXkzlpNbidbQhw15MZ/BQmeitGN7c
9eOmGPStVtoAjWMaAnCXI5qmK3rV9bpq7nMmatLrvopMvIwqUbCLHt1qniQ2KXKaT2mHVwyF1/9b
9rkBSH4YqeL/Qfv62cpYItLfN/L+hWmzvyAwECkfPLOy2liVpO7spQHisOC7xpcqG24wev01WCU5
3fMZjdp6mDLfEWtp2NIlMWMpmZ9pnndsm64W/ccDbmEgTNXMkJGROPy6zyDOKVTIRfw/GOF20Qn9
507XujT0TQNO6i+L2eGrBHk3c7GI52FxP7Q22A/HXyMpSrnLLyK7m2meRWCdXFYPoXgg4VJ/xOQS
2G6tZDPJLIvac+67OCinxm9NmkEKud8AOGG95dDlPB/gd3x6WYC/MhAFvZH04zQUAiWyyYwSq6z3
aDkrbNIux/JLqb9YbSiGEuNJFG1BSxuRNUyD7qjkT0tKWTDAoP5MNtbn9VrwiFebcWZ1MWDBLzES
hn8GYQxAlyYQZuJhNVsjUBvug6+2gChJPzSFFZzFKhRMQBm1IbzuptrNMh/L83snO14DaO5CWrp5
D0RNKOkCsA1Xdzvuvow9k8JK15ex0g7QCq4e7Z49DULDCAk5OrQM8e16FOfWbJfdDjjbViAgdLCZ
+NroweNOcbX3WaFkkyr8ByYLdT+Hp4YoVXD7Yd6G+B4U/m3rfG0xYT31QUE6nm8c8NbNYx/dONvM
/N1ofeRwlMJE6xZkYvMJQjvo2Y6mj2JLuhQthktj9CgvQ5LAuikk+dHBcppJJikdA8Nzn+XFPVa7
TwAbMVcAwqo0L1Z2cXCzaqEV/s01cWOFoaPyq/Huba92pt8wofrTS2Bbqpw8TYn4LYOO0sY17rcG
eXIZHIQQn8bNh9R8UMp5w+9Ucc3r0sbzQLpGiLZn0cswB2H45rucwNEvqQfzNKdklPCiGHKKv7Hz
XDQxED7/zcieaF5z42TuzjEzadcxxH2BGSzFDt/9VxHwWMFKe8LIduP+Nz/lzsZiuTyc7hQ8r1aC
DvrNsuvc5GCpeCYj+SkkOv0/ftuctoJFCe7KplX9l75XyFyOS+gBkeouSxyOpk7ZQHqRZVF5pHSY
Pc9rdTjm9EVPzhLwBWnljhQ2UDnFq64iixOJN8X8DuhPOSlWz8Bb4UX6StjGRTZDrarYLzxEmjZf
oaPOfWRTACAnswoglni8PKSu4E+TuoEjyui3JwZd08pw7ntjneOcGgtc1vzhYhykKpoVgiZlr2j3
av+PPl7n3jhyjaosGNKDTbKEGXGqrdI/AX+I5k7N8Bt+Jh7K5RTVs5a6KGirlsCMmErZxfz21Zjg
xb5FXeBbHIQqxC3rQdizU1q10vQ6DF80mYn2OCas/yKlWbdQ6MyVpGnO0qQyX8IrWSzs78cP4873
Cwgusht2FHLMhl1RGTv43Itrg0OmKXVtgordLA7Nz16E6S8iOXbmQcbqh0Vtvb3fIWLLRlMorn6R
ooSMcfZbZKlFvaobRPJMfkS0a2XS/DcPVsO1ixgz6ZYrJsZfLK2v692oZBEd8tx+7AFMfm3f0hHf
kV7UN0ntf1vf8n1qJZfX09/g+fPIRewIXzBDMesWnTbQ3Bfuxd5XyzgZSvKxNx5ByUISSudkFf19
6tfNFS2aaUbSCTY/CZIUD0jT8D7UkPKTn/1s/6oXgKQOvuRXnlG5x6Nue9gjloSoxBv595IrOyXI
kMVf0EJqadVX1+C4Y2b5sPbgGvNxNKcVcfRoJDtmwS6Cr6txPEO6xjpsJHYzIj7By4TJmcGDNt4d
TOLZeLU8v2sVr6fAEm4KHgalS4dW3OCPH/j2Jhp5FSjerS0WpHykpy/pMz7uJrS3ZZFlrIz/lUjP
VJyXDdF+GkbBJz1o50X+w3SrmUkANdmrdtN4h4n2Z3qc2ehTADR1fI8bUSMczXrMTysnHAsQMsA1
qSU5L3jvXOScEJQ8RnXepVzKcV9RXM65R4LjgwC2wWzgZO/1Gbq8pxSHE4JT4CTgxxhhtmRwM8j6
9OsgZsE7Fr6xSlEUhaoi5RSRXaAWpVWPop2MjCtbe/dREGs8xMKfQqY5TaW7u6/O6H54WdSm9Q8m
9z7nrlOL4LaktS+ExSvzKpsTbkDlnHFKHRMb/C7YiCKjA9bkvb3W9SoSsqnQe/kvy/sRhOpbzFgz
4Mg5XMF5P/j5Dz1tmmW+Thofttbxub+YcnHOw6Xvnn6Qg/N8tvoLN7i5Fq62wHnegkc2bBfG03Vw
+lanQqR5umXbbXnB6xo6P34+PcteAbG+DxNlZcklOt+VjQzKzWGdt4mah/lJLtp221yAzT/AC9hI
n9lyzI/8mqB2SJLtj3mN30u10m2daAIIzBpITZsuSSIc2PMSTCMdha6WLeL3bre6jx+UPPV9seGV
hAOPTNrnlzL8RndmGo+2G0dpWjR2OhTseJVIoqNohq4uqWrGUuI4D9Hp/R9kaTRk5zgCirwToLZM
YXe1NppQkqk99qbh8GkMnmMjUXEjLo4DoL8pcjKKauDE6fanqz3okJ+Njt1/H2NVT5TOnlrZUU++
eCMbdDxwJiO5KQTtRZnNeUXMZY4E3F1/HruW0USNx/b7Dww3EG6sJX3rcXMp1h+l2nXuKob9ngfY
LtGnQ9GLTrGdDXt5AS7TYK411kSGBbYBz0Cd0mCV95dRma1Hcsf0ILdGSsVL8XCxDtC16yvv/k+U
BNZQK9ai4FsTICamg8rRZCOhbmIzlE1tOI4Mo3svg+sG6dfJ+MrPEO6jwOdE5w6nrN2vRbGUbk55
9CJR1IDcPWxaxsNO9WdUDX9flChPBHBEDzLcC5yIxC34BaqMBSxOth1awy5vXKj38H3bf8N5MXnX
TztzQSFFzTvHnEjG+LlyQMx2fr+biRVAKbQOo8EQ6vyleqTVTbE0W7vjtK07Z7NFqkHgJlxrGRGM
CNaDF+3d5H8gq/fOMd87pbgxD2v7hEuJb3qbawrzk0PU9TYLeHlRRp29fUNPYtEtlfPGcdk5oGVd
uJTlF+neZ6FiEPmrIMUp+U8sef6uSiu1xW4ymyxwfrpnYUp3ZT04C7MndAjmbmlVrYm54Egu8+kZ
k0a+1HX4/6gIlyUrTi8lBpuFREg03WR/7+F021iTqMrCSRM8SuwXvpuVyE5UURzCf+8HxwNwzHig
52LdtxVPNq/ogReijOHb2VEKSiLRMcAH7QdqPcJHe2you0dKzuyzvrGrT8Qu4P9pKrRcWThii75R
fW2HMQkbr6b0Jhmzv2UWsh9nqeMDG3yLJSUiGa2t8ev5rrT+epw4+mtCZS1Z+ficHl4kRwNg8XhT
d2/oogiPU1Qcsr6ugbS2Oyw+g65SHF6Ep6jmoIDeongX5E8zT3Y36OZ2xb0ZCKyWdQvDHrkfn0NR
K57JhF26+dQ3ZQ8Dfvdx/PE+6VYs7+9TPsghItp9a+TP+gZ6LJusv0/8xq83FaC62FepkEpCWG0J
jNbjlkKVsF3hyY2kt6BM/GqXAX/aX3j6Nr4G9GAnz1sqwW8YZYabcL9tGaMKO1yb/58X8ZW/MUWd
/VAfWDYb30TTHxEHlT4lA9SsM6yPw8+PbQUdt+CX2tVU48kZ73ShDVx5sQk8gZGZGadvFYR7XIXB
LhukJ9Y4P1BJDRQgmGR5GsAc1v6v10DxGvuLycWpyDePFP+TgR2bJkHn4CfPbdTMXjCd+gVgKL38
lFKOpX8zLeaB5HS4vZgEf+x8oeV2JmDxWYSimoO1rCfQ6rN7ob1guEY8wXHHsvZPCSNIuTBcPYVS
D3S2T6nQakP1bP6diwf6nSdG5IVrRFoJNb3mLQdwMhsXYtWfnTAD3Bxiq0jxajUGMx9hsUrY0Efg
kvgrjtDQvv14Y+H2WrhH1AhBgXwwQKmodd6CjdUkIAdCucq/W3Fr2uGLRy/gfNLoSxpdu4Mtyiol
F7kkEKcDBSepJ2Eonjusf8PMkRPkKrqXrbJeKLY0LJJQW8kNPYPwqhwKYIEDv0JpXl4nsj4ib0zA
/cj9IIZ08TVgRFjz2h8K5TjU6l23MZu8WtF+ZE02wCyDG5dvymIne3SKlDyadrEKRdCDNxd1WqWp
uQ+9TAffs+9QIZdNTMtQ+eWPKnd7kemBP5rrVTS71C012VRE3wDIXqNOLniMuIrXDkzk0EKvf5te
lp5kKBmuYuftZNGsKsD//9DKPvM71aXPcIHUdo44UJcTuush3yIb8SltDP75AXEUUCacOk/Cz71I
R30JGc5seaySi8A6jdQJk5ICh4sBLPkrcfJmoyKxok/R/hzfzaV3ozG+rngnbwvcJ/NWD8DEyKOZ
ZDu3R+8C5M73JECHFn+MQ0Cjj51YGzYvXHUmDEETT6FubFWL5QnzoTQn3WpFit4LMDFZ8BrVXgmK
8QWucBysr+ZEqjGY1ia4Shk+eFVirdv8bDZsbb05ZcXS5uN2sZEwpPmQX1jorGgoGntcQQhOkVpz
zfPxNFMVvEbP39PDkpfUENLqOH+MHDkhgCnonTdBLGj/mLZLGKbgvrxDyIJB1xAQ9HC4Oq4+2vo5
9Ejw1y4nRn+e//hm2+8s8IJ9Uh4x5gblPvVEg8/l/4hs91Y5R/IbajiW+2VPP8FcpD78Z6UKo2Ta
BoJzAtPKP9OOhDHiHlqDEzk0X4HaB5kDa/bqClthxLrAsyZUqAk2Soh26MH3BPmvU/hpZ1wH5GZt
a0GAX2IZT8wQGCaHYE+8TZDoQgEXbmkEgH8DGYEjlbHXbZOJyAs5CezrUayr47xpvTp+iqJb/0OE
JQBEcmEPyN4AO4yJ1DGge/csvWuFiuFAmWDNDp5LD4+fcYyr4fSzbRunN8eezgFgUvE+JwTQ5Stf
q2SSF1okXwGwt/JwEPaf48EDZRYuOb8pnMJBnmxCk46W3n26xFbHkJdl05INtbKHh9FEP2VupcRM
HiZPAKP8L+rpqyd7lZN55pC0+KevEQhVDPIQ/LH8Qg7L6l7Y+1QTqV7qa6Et2J64YeJXYiFWEruh
9gDk8oLF5LNB+4TMfeKeuAdHqnfjvnwEeXS3YeAUK7g2MYpQdkseREndEsJgN3+Z6PUqAlO/ChCi
7TCP3mnveEw+oAickrJk6o7k71thMJdPe0e87V6Eu4txwibme00gwGrTTcsiJJLctZoDc7AIy6pe
+m0ll/XSNbD7/BBxqNRsq+v3xt35zzp08ZEPBN0S5bqEmEd5dtodu/9I28psfRfp1k3rMmt5rMc8
2jO4jsBOY+E6g74IaesTEOTDHF09A6eiTT6qWqEBqoP7Zkfol8Z4xtl3LmdIDfXfzUfB5Ky6CjZQ
O9CXzFN0Yz2hAmWpZoNNbZVymT2xi5H58IeCDXI4wI1lIXjhtymWV1Eo7wKyzx/XCYpQlb+pUtiU
lgRsf/zzOVRIJJDixV1DfNTY1vIjT4nIzpy4pNemIMim1YTTB44OnPsJ2zPBy0Oy03cbrAmBtl2b
ViO+RvejS5IzGTBVhQQFo/aG4do2EPUcx0Nk2CRIx5I31iNpQNOqliZX7tnTPplFvpfADDxfYhEi
dd6eupTPL/QIGijY8e95UXd+6EXUS5h8EkjZT6cx54iv7rvTTvhmkHtcBiQP99Rd2ycwwERmu2v1
hTtXp1Ruhxvt15v1WUQX/RhA8YX2mN/95f4nCSMaMdB9eIL/P/ROyJtYNh1e9MuetsZWummGpcHX
g/a/Tm742AjtZRhrFjW4Zn/cJycMRIr4WgV0MuRRIEedBCxDtfJUNDlqtefdkEmwGDnLIDjQttbh
hbGt1pfO0ze3KcY9RNXnL8HOwn14coZYqNb2EKlTIF2Ze8pzEKdgNfCo7iScvndiHkXLQFHpqkh6
bZ+ZgqZuRDNM8CAQoog6vCR+WzAtolGmHf81y2VxTGLxjqaZz1cBePiqcmiqoIjCTuHmdBuqC2ZS
6fmbc1xeaCGJgJ2NniO8pubWrE2iBLLuOWyILZ+QNYYUYXNXlHXPlW4/FhnhBFD3B8yWKrjE09Rn
5/xXjp6n948vQ9sBxRFecxZiFtxz0WyyR0O1N0rx35g6NL2TStcydDPJ08H7OJjiGY5gW+BxhS/n
4n0xtoJubVY8/MhwT+4+4+qfEO8VMY2DNvlJ1pDp9sqOOkNACXeLXBbE2Y2u3jtwIWv5kAuO5e/w
90YIlnzaVTz0vgs4WuKiygWOyOhwoh/f+TSQY+hJazl8lJwyNzfN4oyF6B9XlYBCKLdo54fTJr5b
Lrd0CF7Epul494+3/qh26OOZHKIv21f4XzM3iYug6lRXUSYR8JDrykBxNJq5yV45MsC0MvbWCqk3
1TTStI7ZJcmLS15G31SnnwwFbLUjNZgRAGGeUudHyMv7kBQvKIjkuNXyJL5FEtCBLkxzDEGFvZ/e
zjf2NCLRzKe2PVDAkkBTYVmlfkQu1vomSzohOsmmorPn9vAhRIwyUzOTbB+GXAbj2RQWt2OjV4I6
ikKoFKGUXyMkF4x4jsTHzYeythApUWk1NVbSip+wuJ7oxb5FSlWSc9eThEb3pMgGFDgOp2+4NSI7
5HCx59bvFUa7zEOfP/4gWgwKmbiBsdV5p7LekAPs/MSEYtAGmKvxbybKn3Y2lp3Vu9V+tagEoz4z
1jeJ6PFUx6BszxLqhFVQzKlLM1OihU+eEJmu8UayGtFFIK4+DhaBC85YUGCCv5uRQXpxsqugy0+5
CVlYcUPIFJA38n7EQmj/gb381qg3lUl2k9Du9oAEEzM8tWVhoKH4JF4GaNa1io8RrEFn8GLEVh1M
h8PiRohaslnKu8IjyBzRl0gq0o3DFJT0+tG8+oq72CmfKcSmaKOe77Q/KYeXKxHamgR3mXtxaq1h
KwvJXQyw7qQNWq9LNEEh/e05bGU6X5hxhch7AS84W+tR5D/nSkC6T01cJ2g5cuMSTH9nIq3JO/0+
gmAk9Pq0LJXhKZQ/KR+/TMDM1FIQtzQK7UZR/CimosIUPkM5IY/acoXgBpwm/0IW+hR1r7R5iaLY
OYEWvhenK7RPYEU/zQTZxe/Aj32n1pQO3/F5Jm+FtZr5mEN754foSMXRFC3OQ6smWZhzf87YLm1W
VdVaNWrgWrc5sVcuOAQUnbeMe/iy+Bfcw5wSBbqVacJ8ORoE4L0JbrnHmIG6T7leIvgZbPY87pW8
dvGxrnZGACtLUUkKcQDDodcxE7gblN2k5QQWKu8e7jwkoZUqeC58Bb4MsceSQDuZgHqhS0psiYz9
NnC+bOH3bbJ5Mw85kJeMjqN2x/GbtwzsQjxz7lkwTZEduy/RIU9YDlweJRqsY1rjDzhqhS625U29
KUYj3G1klXBx7XiUL5iN9j4ns0BnlfweaRQEUomDb0qdqZger07wTHqkNN+xSSN3iDYsmIiyakYQ
oLIpTP2l1qEvO9+NpgFOBaE4+STVwSUmbOui8srrryMA0/7ML8Ppz8ZdYc8dfZJcPzR0kvLiRtly
fGMA0PpY2cE2JIyL6fJjtq7kHCd9DttidT5xYAcZkUsYLKc5kJuhvqYihaF+S554VL7/RTLExUMA
27mCIy0A87WlvRM1o7IiSRSYUE5XwHb2OnJw+xadlwtJjP7O4zo+yJuuQOlCcoK/56WXyXxSlO0n
UZ7iKMlTy3wpn/HwelsGCI5XF/Boc6Tjl9XRt5HL/pRfPoU0iNtzwZjQish9k4hZ4HV9w85e886r
ZKWNg7CVgOZgKPWEEBYJ1wS1LdNMgjgThcxpj52KwtnEiTPSx1iXE0sdznbe1G+88IYdAM0GsEg3
OVLxb9aJ+NUZrcV1181mj75bcIlNEBBQ/N5Xe3HLQk72r8s9qfbAJt7ASqNfsQuMSRD8m/rjmsat
dFYcaleQIXDxCV9k/ckfhNFYNfPQQK9vjxB6n/9HctE4xrd+9jHa2WeCg7V15xtv4w1GMAPyKRdk
DDhXIk9m7WeIl4KrIITw7eaasOkDbiYwTlGll9LMDOuvHGrUvBeZTZYYHOsIo5QpqHDObELnciYf
iPFo8DCt9cupdxcYwQm6DXbNkYME4DMpchSKGPAvMksyF1zj+flC2zNcWcN8ElCVTboeik7i/eWH
wVj66KGNn8/uu+ty7gfGxqjDqzwXKFACTUZq0IcmrSaLsDcnSjhf3TJ6Q/TNs/NGCoshA7LTjLd6
LLJi5+tKZ+c+Rirn72df0a6eqjOynuUjQfsud8sozJa2aqd+UOBvVUymBnJkQnscit2+tlnMRwiS
Uut5qdpUaxbq2sT0hkMn1R7/0LJ0fYMcJFlKkgLEjZAp8bvTK+p6tT70h5MgBQRPdS6co7n3UpTj
lenlwg3WMpa3iRAJL5v/6lqeq1Lr80xG/nBVz5Pupzc7/S5HkTH16WxKAVMQs5/5cghd5wFNkObv
D6VNCXZu+4WtsRgN5C7Tyawwp61CxLapBXIPYcBipH0tSwhbZKRHC4os1OADcCubp9NxeVob9FaV
H6kk2/60wqfO5+2NfmIOkoVIPp7z6YXlQP43Hu87FOlCznPjkPgjiq2SUcaohg8mgfIU7onNJEFl
Ue0nuF8Hg/viGshPN12m0QofMhaTQVNrfSwkmCsjzC4CWK8+XvB1fctJfN/C0+DcI5gi9NcIhoPd
Xia7yt3tUs8tuaO5DVJP1xPUIGT0ywz69kCZISQdOX79164SpT3ZFGCEIy3ONmrdrZX3rSUOE68r
UF9Q99K1+2RMuPTQo6+o+GdGRRELdFkSX/JwnNN0PdItrSfnjofAfOx3xX9Ingp6NEpE1QZGz57M
mF2Mv3MIpu+4j5lrFceLnUX5YuSh8T50Y5AdWS79QrVhFXajLDWn2H9g2wUYDBycZK4R4CmN2HmL
E61Sq32LowlbWvY9964OcJ+izWuEbdpgElOnpUBHajJ4l23kwYFC0mMLe0PSRQnHuUzzxRt9dNP7
LAVQvpiQ8yG9ZUg/eYkMX2XGmQv/2Cxht7JcmeVLbvgw+K6vyg9LAVAjLISskS1ELuvwfiVLQPrQ
2whhlGPTuj3ddiQoBkETnxj20mdCTVzu62Tu7f9Glg0fkkGC5t9GDD5+Ggd09xFYRm8ib1V0AYCw
IgDzgcnBjw/Ggy7Sdmg3mILPfWZqsyXJBkD6jgP6br/jEu1PgF7btv7zChwzXtyExnQbulYo81F/
s7ytDbe+iCmJTkx0h3TPpKUXz2zXJMVFC9L5i/Gcaw/Ac8QktvTu3ObvXESn0iHv+bTuEHFrWYo7
I27Xa/ZmPEWJGNEVHwJhpBPtcGZvqOypguDW1thVZxNpwGRvK518pNgWSN+IBhodk6O5mPxEPu1C
R4R/5rLgsTAEABBPGp83PAZ9mviUfnkTmxMg3Odpv7jO/p+dzodKfcnR9zRY18sGCFhfa/JO5p6i
R930WNsSJ+GDc/jVb4fY6Fun3mIEjRt/VD2DMvF1oc/2ytRvYfsbkmsmKlXGVZaBFVbrZlHdOpW/
22qoSIYfzVAtsAZNzjWz9K+7a2CXHO9eiNs1CrDPitprUG8J8d9DPoXeOeHVX/iHWobtYxEFwSFW
UdMOWwGXyE4uxwZqRiY8cDdOvMambP0ghnF53efgrJmx0ruybykdcmIap140HNKReHklsR7EOBK0
FwsO3NWJqdx2WwCUk1B9Q7W05J3UPWxA6gqHJIphW50z22etX/HmBILwIKGSgqow30puClUqT7OG
+A1bX/EP21+PzLobEJW/eTfIsDZ14NMDIqJxSr5fgXG6FfHsbq+uiGod8FXYPTsT7CBu7/o/aP7S
V/uJj+PW/jayp7mEcDGD6g1S62ToqD6Xhe0lApeGmSbbohY29+/DrBNPL0ILhdtpWvuxxPCKlXQb
PcgZFJOeOGyTQcVg4uLh1yGzP4CTXuKaRilqK9L7bE+c26HaFM/8jUCx4sM3V+3BvS3Tk0xB+P41
wsPXgPLOND4Y6qahjHuDA5DVKZq2pmU82Cjn6Dp5gE93l8BYw+DZAhn28bm42xOIkIMx2xK5EA/8
ggFp6SvJHsNR0ie4aKV91Fw3j7fitceIbBFgCsZXwLXnAZNRhcJjCgv9t1EG9psEjiE6KQ196evC
BsxTms82wiH8AM+ayUVC0TUN6u5jjymQ4J04Gk9WYsqZR8qkh+eMQjCeNoGhPRbdRkiaPl7fENyv
javIxppVzpBOhj4m8bqpcJ6YstVMTaEyVZOGq6LQ/oRvlbiMu0cICuMf1PUMQskc/0fX2LpPI/3L
pMn2X6fv+yJcjg64I+K45wwOjz0IloUOFK1kMwYVQZy2+Itg6gQPv3NQIW7xuJcN4px1vRQefZNv
dplNA/j8JYFTUNA3iFP/xLe3ueaBDfL+CmI7My4AxdH8SHHdzj0im7fuxCf6stdxqxZKjArF5BSq
26InGUqp+qoy9afsgvaoRgagI2RGypr/3hU4A4kX0iVoA4/oG0meXkt4jssbS1wD9y5lxjr3DgoF
Iy7Fz1/thuWGcfh7L/cOO25QlmnBVkXJyf9wayccNO9tSQ0mL0lHXRdu7yL9C5Br057/invkRMO9
IvO25dN2tFVVZdKr7ykHX7D8Sr6/E01wrec+eWAKtOFYH1Z39Z7lQ0Wpw1uHWyuZVBHoECr+mWEH
BJXQuaBx0HhkpMp5tcVegDkfMM8dKpr1C4LnA/SVJX81ylmLHNQjHzSrKguhq8Zqq48+VKjvpdsx
eD//2H6beB4czNPFxu32T23aZ2W8XhKNlhJz23R3NGTTAZHVrOl4APMLxd/jA4xX/JniWV7XJRXC
baKWoTUfDJOWE+1F5Xh8OuvepScELDgfy9lullomT2qsX7i0Lvlmpyw8YVaCXb0guEQ2HzplLh5v
nOJj/uH2MVmCEfzbSOiIGDE3jgKvSNJJLTIwTP2JR/6U6vutj3BMF9K4rt/ZIxvuhvqNDl5gmZFR
QVQzen+6/sgfmQalC424yNT/iKckRRVHk5i9Sy1w5HW9+CwvWhhtr1m+aHymi4mKuLyvyHqVio8t
1F9Eb9v1vGnrkSSZ0ZBeC48HUrmno9hOgmrZ9HYyVv6w71gghg6BnumA3P15MxiwJ9nLESDnsQ8S
tmLozbDA+71oClwhi5T7RpFLTTiIY4wBVdCssfndYk+erWnME297bTFYV0R/m0EsCdFk7UuLh/PL
Uj4VccxvpEAoMl1fkRiQ4jVewOwcR0CS1TDrjPGKvpv0zmh2FHJImyPf0Z8eWgRWUC6zX/EgKFBC
jVwdBr4zKgg2BewzEiGz2dvnF8AMN9yhSvyPJnz4CaNEQVcfGNG1nluQF0kuzqBUatA8t8GS3jOv
eFHTvy0h9FOUNKVnzcwv5Fh1I5V0VPZGsyJU/yHR9v5F8uAKBR/LJnNDHCxSVgBp7m9t2XEtgL6X
3XXxYdgZRfIIMvFi7XyqigYixo5l+S601Nru6end+rdXPuO+3y51sUkMw7QxdoNFbDm0NhFjrR6e
5Hri1uIdJK6hhz0Th2nAbkFObwgD3yPANDUMpkmD9tV31W0Gr6rnttWJq1ZYego23IG3lHIqq2ve
/n5+wPswVoc1CNE9q7ITEOMPvBoXYUnVqG2F/rguYwL5iaoArisIo1WhQDNmE9qwTqeHR02kaTUC
Zbmzbot+Oki045mspW0nf3tuNXFBxWKHoVXB5iFNxAGxnEbMBiZuljvslViUL2Ur92dnlH1pm2je
KIHWo2d5bfbJI1rierrC0rPLl6dJIwGFOjUW2WWlGh4gfLbgHvQpV7D3MGLQyZj8iMY6ZlnOO4jn
MU1ULd1piCnEOBfmA1kJPKhsJKpcT4ZPVxVv+ppu3Auk9hIp3pltpInFLmSpTECNgUHAxJsaPR1Z
UgaMntFcY3cdM4Qk7KbEFalXOarV95GfkeKvxgDagH82t9dg2I2Pxy726NPKmt3TSsXwwUP9wSkN
eDAyUA9DCxoKhR8fyIwggZ7KIZHtdlxhFE1eWW+Je0eVXz73e0s0SXhu6oSP3bmQInI8Z7Fw+2TE
wwMGxfRILkcRd9D05Y8BrWAYNmcBCWlHH3ozdnxAKLoZl6pfQul5AXL/3sSh4PQnx0MNhLSuOQEd
q6qiGlvaI6xTGxA0FkRk7CXZ/LUjukI2+EGJkrAEpcAqYJoX6awUN10I4G9GRXMHqsb3FDcxevGJ
32YTxm/rAiLF5M/RfbcdUbKPhW+bLZvMIQDMWxt0ZyAnFFfcNPrcGKZeY31uKfNi41Er/bLicEIn
fsUhSoZbAJPQDY0fuNUvU69jrpAzEo3b+J4dsa1ZSDpKhRSB/Di1Wot2q2loWZfJKhntZDlmalBd
4YXhpVk9YnL8wWfWBlMKI7srBiddjRfYrNRfc++HkgjV0lhbpvntOVm4HEK7UYXD3MQUHQkOuknj
fqdja3BbF6THhr8v+5yakyeaWUr4e7okwGoMQbFJFUTdFnnhtUrR9WNhb398QHc+yPWS2hrcwTjA
P0IUq7GvdSn+WuM8Nmw+2XMxBAHNwdbSSeecR3U5fYKeFzMd9cFeim2Z2nZjn+U5SYohoaJaw5BC
8NjR+nXrWfAHYjVV26xvlcUjXkzKsrQ6CDMYgNKHeA+3Ak3B3pCEFae7OjHWEFl++bi3i0cgS94X
wA2Zh72wiFu/sQwVGFtvXcrruuN/sqKXSs5LHmT1lreuh6MHiQDbON7Wi8a6qL2TKXXqUsI6CfoP
zyCPcas8gINwEPWv6PP0N/2OKlT1D3jnJtsBReSRNZ9rJ7SesQc21vPfKlBwbAB51pzXqFL1/utw
LWG2NY6Hxf0a3TZ7Sft8xXf4i41qYR/yv4Jc2n0BRwdPqbgFq9gsKLC7oO4JIXdOICAXZwrovJ6Z
7te4hYkK9C+J2b3XErddGdSEdrWPJcV81KSt2lAUhDoCuBCxqguCYV/hqNVskdmUV9+6nBsJ/4eZ
PI2ACp+U3YcPOjE9ggME4ys0BI517fjqWMF35uvOAfZVDAo1QCV6Tlk0qjrhFifaSm7gacJZZtxx
9HvIlKasvr1keZAh1ku+RRnrMWC9j7D/daWQdRrgnHFMBS+o06y0s9pQ7nZLF4u8CQd6CxYX91cc
dJMkzqT1b3nOzB7kHf0xvhE1OwMnOL2uB22XAJoCfIqjvh5dNuvnvem+U4HCe2ZJhq8AFjEBGLnd
wvGwcq8p8GVbdKyNdNxXQld2N1okFoJcfKSfzDRc9g+IZ1XL/V3S8Vjwx0MSqj5oSqVf/0Ak1IWK
33rvF0VIxmm1YQVM92TjLZbVky+gLQKks/b1O+BrB6U6riv1hci4TyCSpGnt4Og10JUyNdExDVrj
ekN3O9yue5APz5222bGbN7u1dJ/KjvU1SGVf90ngBeSsFwxfiylU8b3X94FpR7VsxA7AmwlXIGMS
+34pVqHhT0SaSD7XQ5V7S8/geCYsxFOW8HoE6oqQVQEaFCLXQame+Wp1lwhEJoauZf/N4pRSXVD1
dp4ObQ6Ww1tWNcx5VVZbm5czFHydtqQA+aXfCWLswj7Zvf90+tDaLgCQhzh2zheuPdgDvm/liPNH
4loI688ozow+K3Vs+1CRcXipMOmNoSR4ryoTJfIE3c+GvjUf3rD0bBhpCPTZL0eiq/sRfQCvLudb
OWVehbK5jJqrFX7ifPT62/8fvH7Wz08Q1a4T8jD9Gmg+2y/8KrJcq/XuZl8xQNqbZASzACiVx/p4
P7ofYrz4b7My4nHu8pwNUGleUozw6QSHIqbIXH8W77LIXF6UjS+eM+EICZBmxDZM3aanDosSpEzs
kWjohIp1t0RqZooKxGUTS4Ekj66BZRcm//Jv3iDhakMaqmZ6AgQDg+4cE7LdbCZJdenZWhHPcPvQ
svvtu5jdYsNwpg7zq+EiymUNV30qsJ1TFLXSyxjScmp2lS62rvuAFbU1+P4njBUkHUbziR6IVP/N
FFbA6Pvns5jFQ4mK1UsbVZGdrt05M2tnZvosMlWsmBLiPR+waWGiH9c+b78JI5F13XSpHO4uDOKs
XeJyxmh1PvC+1qry7HWunbCmFeQferuWbyvsAJujnksNFoW24s/QiXKbKqKfv00b8SHR2PxD6K4S
qm4dCIsJDOoxJvCp6gE6OCcBZMdMtvKcG4OEl3H0AgYGzlGY/N2Tef6UPLKXx1sCOI+ranzwb1a2
40+ROqT7PheBfVK8dFhgaPdxdojjQoiwB16bZXB5JtyAQUspVIIc9CJ4+shCf608c7DapFR+6FFv
m1TqeVn6BKVFb7IWmu8NEeR/2b3pIzQwnv6Ppsm/quZDgBwzpHWrWE6dCdRFun0BnmTJdAlDeu1z
7LYuIJyUo5mSkGjFamaMy8X6nr/k7+5mlPMRTj2O6Ub6GBSX3bqZUWEZBlM5JAS4VgguxRkZYSH3
UvPLNfbQ9m3zeVrTbI6DrOchYNUbDs/7XA6B7VSxsTUpho47IepaMFyo1F+rgbip1l9U2c6GRTmO
02T9keddj5+eRe9MHovcwbwgMqXki0KS9VoLS8dGWESS9gnVTuK6odpjM8RR8i5wo/nxSar1GSzt
zi1xM0rI0I4gAgwwTnNpdUGEi4vgyKoU25sccrBuKl2IqioDZWQ1nL8Hfr5CKNkyXxMg2S1SMPxk
oS4OKFp9Rq48Zpxnx5c9Bj3loHVnOyH1IWBhJQ2wXPZMz8eEUxcp9dkMogMJ4qJdYrqFnCN43YBS
fphHPvhZm1xfWq04RaCSH3Uzw9FMGtiwE1w9J5d1Dt6gQKqS68UVN4BIM+NpzGd9DtuvXWSniZnC
Eol8vPeUhjgEjEhsu/H/x5BHGwL9PQYAknZgjIf4ga7vwBcynrCL+A67KAh/JMAiflxNwxgl1KKj
L93tMu/DfzcLCT+G/jukqNfB+OgIgUMo3uOCbqw53nhj3htmqjTpNf5sf+CMSLodTZlFR9sIopoi
wKA1yABrEK41VgAgXGV+81gOZpMlyms9gEVX6PrED3igmwihFFqGyL6gQlhNOaAbbHAxNPxoLPtt
NGEp7vq2POIM211Im6NBmufG+xQrEWYn41G+WnihK0T4n4xe9S6QlN4lnsCDBlzo/eee94drH/bQ
TznQLrB5kOH73yjv+qKIbb52mFX1Jf7a5f8F8ivlafdI+p501IbzcagANBqPm6BVcd+g0C+qxGC5
P+HC2FrEgeCuTpaxy2UfZog1Yl+JAmeU1zZ9LRTZHkJ/E/T0T4x+pjKvIfqkooUggrngnGixInSb
mTNISVWk8gctsM2jyZxWnWNdmKH7CQ9QnOiTDQ7LdurnbuujnvQPuG2iztNX/TcS2HVyR0e2u85p
XEXvukY6AjNL50/1QsJo/wNzflsRFlbtqim7GuJekCAQYwSrbK2TmnqzkEXiLnrq1uL4NV1mjeS3
vW8XglGiHign6lQDFXPzJwHmmhadf1BImvmlPa2wRicXw8hv8z8nFd1ERHj0NqZ3e4x8DcwPXq1a
dmTO0m+aRKXW1V+Z51j+baxfg68oV/nugSRaOsJo52/g+V8x0dZ14d1QAtv3x/E1MrhyxZLIG19H
uvf7JF7ZMZfn+3W5PZhK+pRcwOiUu9YQN84S/iUuXlmXaeBxUEgKOzMFWiJdtlRbkLqX2BjpIpjI
FohitlssCEg5zHbuuTsE55V+2Zyi57LbQYqdnmMHzgGXBJ+WGBOPLwpqRdM0V0vfAIYE8HfHwgX+
BSM3CTpY8zvSwKAdV4k2fHMkkI+MmUxNp1VMQBgduIaQ2pnlLxPxkkY13DgMyuK2ki9fSYCEiwnJ
r1XwM4hkRgVVOBZgOWhARateb78dOqgTgCpmnzLoTwIPcYv9hU9AWJzTIAKOT7/szxrQZDX5W+lK
So/YeOXkyUsgHVvtUam6kxgU1V68o8xvYhkfXR3vMYBVrc9I9nKBvog8KEEXOWBNk3wlj3katqow
2ew7gl7+zU9W0nnL8ZdqnwqAkosy/pvsMhiDRCw089dN/UaNlCbHzlYoTJeSOgOw55zW1NtzJxLn
7NVX5Ab6No9qyVncZW6hGEsFO0kDRMyrxwIBc3fnjVkHlnjeFpwXGhNE2QeS4EtTnXI/KsvZHmP8
wFR41Vlgw2uamdgOHvpnjqwVpR2Ax5mjgNnVq7PnGEZmutyyushFavQL94+zzPem6x90QNhPigsZ
O8ewolCaCOu2bk6cSwm+eV7gJkF2K1Vhulcm44SfR9/bvGsxfYa+cn7kMUdW2v6ItIwnEj6yCZiy
g/AO3XADG4gQ+Lc5KmhfFYXUmmrdK5pUDXAbAF7sJsRjCekoxQXpjAC1Ar7JWpD0pM5AK+pAbYZi
bfyjcQfrw47llzulrOeuL6Q91IYHtor5BlU0fKhoadQ6rMWlMI4umF9RrjrKxfth7G4nDpdrGMHN
PCIuHrUP7pB/3bZzvmOz7r8aBdddBZc3jRHnsm9CSOrx/1zyJH4kZrsXQQIGSQj519cFeByUoryG
BVKkRazD68wjhYOaGPfbapjIDCxGFvEWVSWunv/NpPHhCrr0p2j7PAj0638qTymiFWefREDZYZG2
TGjviNKUN2dO5XVxX9eZlgm/zW3LpVW9bT26J+zUaKA3qFHcSCY53n2t76kcKNBDKlLMMPc0smIY
3YnHzy+efrjh3d8ZUX023tJmFO2NcFDapYxHUwjLsrJADtA1Kqvx+OWeDIp4tmIoSnRsHvHRyEWR
VrAlmSW/bUeIq9Xod86wzlviLCevwqPfK4lpHZS9aQq1d8ibOq6Emqg5v7wgBcBpw14aBBZt9SQq
comUKikQw6JsvWD1RKim3si7syVOaWGhI5Se6WAn1JxO2G7H0uV0RvjuSjLhi0lqmnowWVvs7wk/
3HgNqGjzdPSM8AnQnu4DCEAfY3ew9kIY+Nq3IZ54S+On8D1108ee5VX/xl63MmtP4NG9y9HfDMxG
OJcjS1lby4gReSzCTwFSTF8zuGSwxeAc1rcACgksVE3pSIrXA70Kdw1P6NMWnO6SeQS68jTHy4lH
RDmrkEAEv1DNH/keKmwoAzPyGtz1rbamc+iPDyvTxiQV7ulNSz+FGcnFaSc8NJbTBsu2xt/Y13BJ
NM0v+pbD8nW+JELHEwSbPq94IKxUxlx06Iv2e6jxI/b5UmkTDReaXbEtHsQkqwI7KwcimudwPyNI
m4+5VljH6eZ0MrXw5HihMK4IEiqi5gSUp6o1x893aOHlssVku2WFhjqgd9rqnh9mmKng/nZtsgPh
AjSgxMk5nVLUdtHE/65BGtmr7SCt6Jvk+NvBTibripoIwogsEBYcVUwppzT3xbueLO8RCTL4W8yp
JIaKEdRdRs3aUDwMICv/DrHAMB1qHN3FYi8Ysh8w9r+R9j0tf2tDPFrR/38fhq3qqkQEsGE3bNEr
6afg2ZseCBoYigithHVgSwqN83GItALS9RRzgvRP1Wj+YGJ9ADzKVtFwnt9DdWN9lKxlwvFyA8d+
//PJBV/T0lQTt8y3Tup/Ug6KMQdeBW9nlBjgZF718+WHB6e72UbOU0NEPrHA8DpxcnYRSPGQlQTw
8g4uNXbRlw2u51J5STprOMhUE+eZZN6VKURXR71qLYaCvDsI9fhHwz9dmPHnXTEUXkO8SAD9UXZQ
FTjcfR0GUc2EG3UxUdYi74t1Vkq6YA/LG7HFzG9FIDH+BP5v6SQcyNldrEL84jPa1kC3GY4z5eS8
WJ23wArgtiAakSbcbE5VX5RSZgT1be1zjVG85t6bGBNZEVLX3AeP/wPNybS3Iw/JHyXo6ICIG7BK
wHvkqgDXKm+GvtNkkf3t+cNF2YRQsCJjJsrPIlAg7pcIyttWHIc9J9HaZX+UPp0vJx3mZ5GIp7+1
Ih0UwRFnhJBTm1QMQeS1Hgxjh4Xk3xaSymaNWk3ByOfUb0SKBr/pLT7YvHHw+yJKcuHwqjjAFnqB
CsnzZmKcQ0fzrw5nv2SYeo1Ex3oCtP/c/WpmEkvyP3pHDaaulbxXnMSns6O9+n6kGXfKGXKoEZ+N
uAfR0Kj3FeLA7Q7ZIRZNxxigIMCabA4fA/ArMfUm4dXPP5IjT48Q/UluRxSXIBuCMNW9IpUtZ/9E
bzmrAU/Eq7DVEfmqCzhv76rIjBgQ6r2o4pR4JF32jksRE5HwQ/HUNQjaMrVbc40q5DhxYWRBFeyS
93xriQ46OKhSdcTrrPLSkfW660VI+t4Igdmq/qPxhJKlGBq268KBo/HGsmqDN5Uye4bfOrc9fjV/
fsOabEwbdzwmuMY0kb1fzt/zS6A1mpdJi35ZvXcKwBxBp6uicPsQqHmMXtwoYxyu1dvfngJreDxT
GuVbYD28JINzcYi5R89hQwSST4WwBGqoc76wNHu8xRXpPtkjloZV8y8ElP165mnxKt0/hqehhd7F
p+QBzbHo4y4ElQ/vodXWFET58U+yq4hDnX+GTNE6CqHUWq+PKMs6sR0mFCB5Rl2PGW6pYq/KKi7y
4UKT+Aoaw3vAxA+if0BvFpIP0YhAG2bABHCSnNoKFUPcvDiXkITKZtQq6rCdj3+jUpWc/lWugszj
9j5YDboJRn8dAd0M3Krv7/6p/r7/EFvzjVJmbb56Uf4Z2sIhw+sLYEucSL9c9zLKhSCyfecdDcap
p7nk63udpp/fdybFl+HkmIRL43U65gAOc07igfgwjqIkEoKHrfG4dHr4hYXIghLIVYYhzJgcV55o
1g4jllOnTSgAhs51PGr6/3P4R2aAH/yY793pjEw9z+K86k41nwEd8u156I9+do6lYAjUvPt4+aQn
3UHsUYkyI9Cc9Jwt+DgaFf7jE8nOw358fCLjM2cqDTzVQsJZIXqvrqthIbnhm1Dim7HvvnDAg0fw
ZVIVaC8g0ygHm7o9efd2g9A1EB4N2CtKAmz373GXlUIh1+8t3Ice+m6pVUQp3LV4U9NuYcSvqY5J
v8YMnuNO10+0+2M3yURAnikPIi6DwxSxQLgceOlzkTiE1O8VYjKoGkXA18uKo2TxnIGWTE//S937
YbOoXk8e1NesvoXw/4kObiGFJg5EteHB4gYa16sUeg/1SZajUf+C3VSd17ebJ/xm3H680I7Cntik
9cso0X1U1QBRss8JhjtN2bu+CEl/V0HR0bjzP6OA3Eb/nh5Eq7Vw2mdIeD6QqjDehtsV3rI0rPKX
6t4/+JzNNlNwJbXgcdyq0//i5iGPI1kNT7ViLZE0fOD89nOiRLCB7GkaOxmSydzZrZO5pb+0Io4V
frFTxVO2C61dP7YSgdlDFwavd6tJr7RUiUj13bv3YFJvYBsC0IM34hZ7EoavOlLMFlblCisRXWSf
1ka5XJijtIezQQhF5Mi48lglqNklzQVC+rxBzfKVIELrxCEpI4A6Py5o4NMWuzVe3sxA/EJrd9Bq
2JnDAYnkD6vShUCnvAxM44VRy11cemFdDNcxCqsH4wsc3zV0jDBA2Xftzx1+hmPYNjTri0AGwfOZ
HC96wFMMUvLlyUq971X/o2TsWfVk2iS0zv3BZT/JqHKBymLFD4nWCBK8jgMhOC/o8OZX9s9zL0Ee
YU64gCU2U46Kjr0tnvg+OCz7TpaD+c1anI2jvI6PJklWUoTyN917v1jd7EGieBKXqr3mOwwmFVMV
QslzK8oABc6q7bVbccE6M0OYCnV2TL0AVY1HN8C+qsv/l8TJbIUIS7DEG2It/O+vQAh5G/vYMgNU
e0WogwhGJ5GNy1lpPIC3gYj5i18L5U/e1MkNZ7AXunn/VFYTU6VkKgQ+4ZM4pBU9mkjWZVIx27Eb
i56xZOI5Yp73/q1MA66bEribisAcCSENvG8KX/IO9IQaS1Ngt/0yFGvAPxGjsJV2kaeyG605OcrS
avq/c30N1mGUk9Ro0STVUWriaMSLCm5qdzAV70eHW2vu3AKEVrpDt3VPuBxHVL95ocZOFd2uloT/
ZpWNK/MLjh26VncVCFGDnGGqYegZGHq+2dx5hE/clQSUS0g/3ih0n3S+brZWtvpx43lHN3UCLPER
Z847UVKBz5gSXP+vGE23GUkKCO8L+Sru2gMAeIMPA0hupj0zHyxPNaqcKNxTBBd9BRCjbj223Fue
fINvbp2zMxjL9gvdrFLrZmJoicuGTe3uUx6Pbrg9kT+FuTYssuQ9K/Rp5OgXTCog8pyzcfDVUREN
BeomkSxNM3NwPhh5UhnVfSrXrBlXUktC3fWuweisdiWSDi5TOlqSEz0vB3O+Z6Yiem+O8A/y7Dgo
zKwp8I/ymmtTqtP+H99Lk7GXzfXIf63U4rHeMIxBqF+2SneO5MSR7/Wnzp4h0PxS7TfTblxDIBc3
heRtIPn+MigNy6c9yT4pjvBeAjkPJo/2eWGGFYmRvD7TxmKfcxjN9aX1TnfxdHijNoGKVxhVRYIt
hymV/cDfUAN+71zdXu2shXIpZ/ft1+lRARaTsxIKnwvYhxonLGSOtZiRkLphAHYYCvs3OXUtD7p4
KoeomN1amfzETCKYUXBZ2i+eF3lN5n2yUhcMTkhtI/HmkrwAgk0W/SKipcvyMVbDHHAtTmYE/l19
avlUvb6ue0gIJ+PIfutTVfUG472np4a93lHTnHbvhG6dQiNtQR6+hy/7UKotmLDPFlRQykJgTsyt
6UUSCu6O/J9DSlE/DygAEIGvFOgOgKIMn4jucM/CVEn6gpBKYiBd8ImkCDt3ZuNmnU1M1I0WX1HG
7eSqJkHxp9CCymadK4XIUto2RzVBwHZbOjEK6XM+hbdm+eE/+HCMhP6XE7D8cHUalKHNYYmO9e/j
YREmX84Twgs0PcN8uVGy/WRkSl7T4ghRMskPMv4bOLtyyIsL/qa8paZ8+WBItPE4XYAINNEyXLkn
1LI9z9hJHYe4Pdnh43/GtGhKcLL038zo23YtnvUzWU7zIUR89arbz9Ze8n2tj0/BlcPJp9k4ZLza
FDBgsiO0Tz3LeFDVr4moimtVi634gM8YM1+DCQqg4HdEK++xnweipYz81b/SvUUtfrdg9wOHWpLg
cKQUvFG6JxnFr6j68Unel6Nf/v8wue5yFwGsl5KcaHFKFk5jGiXJcNExMxhIy3t858X+9WyZoccu
4hmAac9AQTtVSrd5l3Gd3OkNcsFuSZzDUKeBozUZ5jwjKXUwrefj3h2qmBx1oALQ3RC08+CPtDx/
wSXzMcZFG4NGQ0bmwP9kqVWib/4Fbz37WGXMOEgXL0GIZIotejqYXsptvR7oPWqN2zay4pySFBHk
ZUhnwPvvE/3je0BEu8Ape+GZKKclj4AW568nHds+pg5jiOC9TN3e86TEP4U97hreXyx6sEa/xW7y
BFmsDsF9zUDRJBck2zVHr1mmAUklMx0UzLsyhMKhq8Y61YFzvY7En3mvNMVYY0gqKd0ZXWYDIuKH
eLC2VjabOp6ebIypeyxhN0wRdGqCRpxovk7dyGtBVN9koyB7Y7/J48zja6YG8vaPq9okJ8Po+KQW
aN6UgVZI6cM6Cqkk01XrfTglt172QM0UrSTA343Yiw9LiZSL/ax01UhRxv3h7jSSZMlaQDsfK/G/
Top4hXU+rFcHUZwa3Z+ptdHPlliEoXO9GuKxG15E4GotwWvhUz9xMhOClLOAjL/eHvfLJnyB/Rao
ZoF9xBP60Obwc8+KJH8w2pY6KCX+FX8Dxce+oiCDx8fdPulPswl8rbvzaneernECyRQYwntQuI7W
u+UlqlY8fk52LVjk3vgtPeu9DfHVdUQnI0vcfTb1ohmOdF18XWcH2rQAoI4qCgS+7y1g+UVkgdZG
nxxZBKOttGrgU9JR/ubt+5z9GRtd/s2RR4z9lwEI5mNPj8opXtBAczZ1lU7Xr+GOdFf6tpn9Jik5
tP7NO+swAVxw6MtNVPDhHmkJxugNCf/vciWe3a3FykC0EJxWWybJYyLaPtTJJCxYQD/IhUFyFx40
t+EwAx4rAKhnR2vy8/ZCkSCnQBM35d0Rc0HajhIZh39pC9RxxsTbC/DriR0h9BrjKCIzcDuPPufO
cN00sl3XT9aRLK2wzMHW1OORbp5MleiYXSv8NgzWQwAp0FPCry5kT894ntBJ4RsCfhGg7X+LCfy9
n2RovGIY+jiHFTNE1SNb6lFGiAmeEQ0xhZeAhL6AMs/YI66wzCrLj/xwHQFQsKYBZZGvVV+C7Fae
0XAT0ceFtLO4yyF7hiy9sqx9GW1Vj7VGlJV+MjY+h98zRzZkkWg+eJSw/9cu2iic4HTrYiIHKCNJ
vIsHLwvNG3YVi0SSo3c8Ukil1ZVi7medxT+7QG4aBlH62/CBMe3uZ2R3HOqc1NKZFqA8xtpuvGJu
GVzkBZyFriY6TmFjYowWnuw5pgxFKOlp+JD0cj321oA0pj+3GXxYvkD5dMvAm3CLXIrDdxaofhGX
lPA0Aqs28fdRKwC73Mps+jbAx+0IopIVQiXRKZ9lHzGBuZGhC4QT4yGLgxgikE1xQtZOJcI7mQ2z
+ZoJ7zkyHbnC3ynRHNGdwEpHEwJf16tMXWhK9QB2F/HmR0r8eDoZhYgIhXAju1ZDq0rd1X4+Lb77
BqPdzHqADIsYc+xYmPokV6LQE5V1wpCK4ExxnyW2aZdUJruxZu9hAeWL3Pd5zKWnkZVZJnXdBONo
SqIjxzlQrywm2S8t0LzhOdGBP+m7uhSVis3TDbuqlg+cpOVpA/2dyRhv65Hb3XmSDgw7EppkLBya
BqcUEHqvRkQ53CNJaIxfoAio6jmj5jwk8+xFVWsKYjdCmprzEnXfYKkt+CY0+brxcsThoaB4lmQT
TYRET0JCKIG+yEtwzRCxEzh1fkAVe4wJoWwKGwumYHRL8sIM0d5KML+pBKOKHCKgN2iJ7XHDC0tT
PjfG7Bz/GE8dIWZbbK7UHac5SjxwAyPJLCGtUeziL1p6zAFSJayP5O5gdVGy24jSpoCfryO1XzGM
rVqN8CoV5QMlEk+mf3ADT36gJpw7MnoqVp9JAjt1hWPlCf5eiM84O/ucP8NTi54Wu6eSUlHIW2Rq
doDDHODTnLxjNB1DlpPDFuRkuahhup7Ga3A24lEX5NLXWpAKSBWQs4X8wptadB6/TNvLgGdavmt/
2fE3jZOJDd0fLiVjj2HL7u+ATNp265zEp/iymOzTrFY+LWbj94eqJuMiyWgS9xIYFOOoLM4v7ATW
hosscmCSnBcxPxDyrBe8OBitAy4+pbElZdGRq73eD/afNoLNrJFh/Gd17aSf4LrCTegTOgU+RZoe
z7Pg1r/x89sJSMpNb7cLIEMiE56NRAAfNpCGzxwShv8tkD1RNzfjFBF9rV+zvgYU3Oit2ZCFPPnM
9sDARnId7KCenHyWWgF9T3UM1tBqTFMKYGj+lOzUSRFI6fIouLu6cmERBufxbvg4FY+VwCUPCVPG
fSvAA08RuP5Hgsc+avCCGbL9+aolyp4Q7Ssi2kQalb4oEgL6qfpZQGiLuA1CQSpGMPNbgSio0A50
IVK0MzLZPg+kTxq6ynVxQDgVw/3+jEspD0wB77c1d3oFMIh/Qavugu9wHpHfmFe0XRcYCs9msP8/
x/ZytpjhJzsmbfuM/UUn2PS0zE/O1L6GZonu0CFEwX/mGhRVFKlIEOY9/wY78+4bIwgvL3b130Gm
TBufepBV6W5DdCCZB/7qsjA2OcH3ku64wnt/mu2h7ItnQAW8Vvc4xNeKBTm6IsKagmkTFJXWZjjc
Ivu76ycRHQRud0x6p1/Gs8j8eGFlULkcxqeBT+cEFd6HP7LAvNImBLazUPiZKtr9A/S9oaA4u2Eg
JIMVGcOvQrsnUfOShCwZhGhO+Yw+Ls1S3JryBAadqtbISY70ur7GeYrfkKgXpj46v1BC0vTbr8Tb
RYHBISwzYyZf78eei8c9vW02HJ6mTCp1iDXPxOrAfWxrFelrV7dVe/EiCJmLn3a+I4MStF4hICJU
LpHBxBWWYYet1tNaD1SXPHzty82O9XMGatD3Or+xWW7hampgqL7W1DwQUj8w+eGF+XvSxRF4ET1g
nXGoxfzyUWYYoGykijm+t1YE6KBCznB4ATvK72fi9SGEH/awFTFO85i0bJw3uooFsQUycnUxveOY
IR/ldAFcO6+WWS8daBSN2jAejPTU+I5j9q/X062PNicDWR1ExXM5HpqEiQkHPjmLU8LmAARiFeHb
pBSbPQs/vhv1yjCaJu3XDWjcgqhK8Aqfq6jkKIolIPL2lDwrKmBlS39IueUnOVP5tJ/CgDZHvX3N
KzT/bKoqJuertwvTI2TC6QWv6NoQdqaeHtNB0Nr2y/tNoYOuKrOq/zVhM/4lAacpx/DZoPlKlnKT
L9DnhCdv8a09/V31ncfyfIhukSwkI8vV3X4fmX46nsOsXn8gk2di8PwrWck9Oz34tn+rTeHhcuFK
M1qSpV04LBNIP52fDmCBw3zFyREAVrDqagwxEEBnBq+uiLcYi5LHKwHRn10+QtaDiBV6pjnNKhFC
eECTVI2QQW46GeksTUnsE8YNWsfYYCiRNNzi1fOpeFsYO09B2H0306kKz7i6J6QiSae6/9HN0Je/
l7OkUpAYPR8hR660tWwFOrvTqua05sC5onztB8pH+LpGBsLwXvMOcZlY0cUS6wRfRvXqPmsfUGVg
eSGH/PoqaZXe8va4/pI4BIfaxGmeLhWPjFSDX2wlOLIR9G/NLO0+Az6/g5D6K9fLsjOZ2FSOagKI
EjY50I6VdlKLrWDaT5/f6Doj7SN1PZBuYPauxiIfn9C6lbOfnPe4AhieHnU2XjyKk8xnRWM7JICJ
AkxtM0ft408mkNKCWCruK++gQ9EPIf+fz8XWqNsOqiG4la3krAUWCP2V/O3xvU+QEktZYf37JQcv
v6Fynx3gytUVOXOrJDaET11wrDdBXha9b/09L9Z06e8a5V1/u6dO81p7jnfgxOtrS0mOJ1IrYRk1
Zv8zqnf5ZEzu4L92QbdDd8ZzLNw89WsLmX5XJKvraV1AGH8fek12eJyMJ65vXsZ0Nf5PIZQktpCn
gFNVbF+sAbiaEOIeS/ju0hwwAJDTy9Nf88Pj8AytTaJCuong+Lo94DT4I5bx+yL6gzgU3oCwICed
DCDFdZ4Ns+m9KyZxGOyhv0wOHYshaJ/GFkkkqkAuQKky0J27NIYHv8FlWDePKIu4JsZ50Thhxtcp
txqtWIcdF0mDbRfZq+h8re2SvEP3bSD4z4LMoxqXsVJwqpMwXyCo0v3OUBhgfXZCGYb2TrSxnXzL
feuITJA/DAiI1Z4VCnbC+C/sZHM8jy+31VwoMBkCso/7FhcAjHJdO0czkoq/Zb+4/OSg+z3Ru9k6
2e3gziMUj5yTLNwnk5TkQTEumrFkSWWSCSEqqvwlgQ11ZwKOmXh2+wlxM6mfoPwMhkv45OuDwxpV
Xa76vwjlWeK396ZLHZ217m6vWgsomsWhJ2+T/NrBnP9uX4Fs/EYmFGiqD+z3DQBL+WwdnHa+J6jM
hCN5UtzpF86rz3lYVGnpm4nBGdZI7C3xuG7nE0WTTGaG+rkNjGBBqmu+aOY9smDLPjFmNQ/11bbL
yKvL1yZeHy1J1d18C3tNTkxo9r++4TOnyd37ldLmprS+6PB+Nk6xQyiNMrPstSbe4jM2/1p7U3B6
6VXyLbOTKSU0HX3/5vS4wzIciSlsjRfXf1aA91IgZTgEUhzddA/FLWf0G68JcqRjunpkAuX6iCXZ
Z0ueiTetUOXvz/d1qnhSkJRxpfy/ywySdUHq++vzi1a2W2H6804vdqRVz8Rm9TO3FyU9MU4tZExC
XgaIuox/9WYxEhBZ7UgK9cg2shfgyIndpFUoKegTKvdg3Pu93qqeR/SxVg/CoB9dR/1tXjmBjkiM
apcCfNdrOncx60rrSCahWUuZJV9Fm4NpBUVphFc5rMDPQK0yOFoLOcxVRTHZjm4Im5EXraSxuirx
WRN+5MfgMVtUjTFkjxi/Ic3hBOs69GobeReIQXZKQU/AClKIftZJgxl+YF9EcW79MCpAIh+UTT8p
R4lHG1LhKO9mK1ZooQtS/T70SsWbT3MzLvYGZzz5ROcAqPSVv4zKnIZKfwitJctcmld04yHMQprm
QYLeaLTci5P3jLIpkYfhdv388a7++jAU3MNF7d6NOhzW9K9JbXrHZHJVBtS9HqCrOM9i2Y1OVQJX
OmjQzumz0bm5pQNCjTMW6XfpHf9wLq8WI86C2Nh9nzYFfsofWnudA+9PoPQp1r+G0EcFw6RU2eT5
7WWKzOcMnvxDAFEmQ72M2ZXFODe9XiZfmd8E7gJTWy/rD3v0swPbco9TLeg7QVz3E7yw3sRSXfCY
cpfLpv59jc7nM7pjfgCtVQlqlYztQnZVFjK3lFrKYrLHjWyqweiTjDwcbnTNxkaoPW1bkDCmTsjg
tcLARPtBod/evSHE3O7Hgjai3F+Xlm2cbsLIF0HDcugd9esCkz5h9kKcRFViqCNN+EkiW62lZzE2
SJ3RHqQra1N2I5PgrLHoKRmALjpWcBsF/6MyK9+0PJAtw1RlanL/pL7qjb5xn2Domank+YelxuP1
ergYctmNckczCCxj12gFjfaRTUIsaksVgA07iBJfr9+cpWTg4Jwh4ZR3Pe2/qXzqbyvZUpf2Zs1a
aY/I7psECP9zUBICkyDdlZS/OZOQHDGAdHMp+EVev8AOIu8IXEfftcrK1GnbZmr7xsnxC5iusaF5
Jhhf7mI6FFkNCXkHhEqO5Bjl91EfpdJwU31o9YKCDKm98AW6aRYoIcXOX3Xq46lR/+o1wcbRRjWH
j4w6+mdxDovt1Yi5QJQjGzL7/vuaDEOChS3zMwy7GreIPEHWqhyuX3IZdexO/0RL2Mcn4jT3SmCW
LnR3VBCPzShrtEOFo1z4eDt5YdMJK2fphHYDfZTKSyQjxdy/1KSrp2YRN6dXkgJKRxZvxD2mzNeB
JDaiTZcP1m8LnWHRke+GSli0ui7guTn+6ygGaES+o/8xqnR7jMW93PR/FXVVoiKMvig1vlkMBlPf
GShk+GcCtZNUixWr6s8o8ZoTyegmdWlRUGovvxViOoFhH2b/CnJP2j6u+QwTL61yMbV9yHEwEvEo
Jwbds0FXx0rqNRRsILQsgL0j6Y8jVg+RPz625MuBfe9+m3uC5EpB5X6t00FB8QwLA2llVJ1PLP4G
MDIHf4o2dndx1R5w3DfvrhvP7r1E35Zh1CvQMtZDoabtcr8Wbz+oVeXrVKhIHoek/RNBe3UnzeDw
pcJ+IaKhfh66p2hVWEtXNj7FVkEKjMpm+ia+Noqmb99oeoud5rPDMnDEJsr8EUln5W1JGvsd9R72
bXl1XA66f9IEv7f59H3fmpRv8aLL3TSenPn3+0EC9f/h97DEZKmAy+rM7OITa9gH4v/e3WJYeiSI
tp/t3N2zxiYuYQ2Ed+4iByCE8Xx6a9nj/i9e3KfOthYCok4jRZc3DMwAwu8owpEd2qROqzYeRxd7
gLq3dP0xuku3ChNPu4IB0sF6RJjzgwZ3Bcr7jTmJMSpAwJIQxI6oaCZCtXJjNNzy7KJ78Lc67H0H
oFZTjmDUqL9/Xo30KLKliQHe6coMsSItoGHCFGArZk3DjGAXfa+FMRSr9R6/guMrfgC65es6a/SV
+V6EpJjJiZNJ2D9AeO+SFJzrQTn0tPQG5mGwnj3pnAETiAZGZDXLngy5NXMgnDW1LXNMgV3Roddq
+iFWQzFDdLnkNMmFRW4GnkWUeugNIgiIXsZfNT5OdcQONOhrYZfq4GWaHhetMMpQR7RDreucESMn
/4AX5aU4vc5V6KqpK555izKthGFofcYknTeT3R5nnlcEO9r2k0shl//g0LDCMMNZHAoYRHE3stpJ
3O+IB5geIXiEGd6dtj5M3hYdY3xeIDPNeFkC9Fy9qSeGZ0WL7TR5Gze3lVgpU5o+2pWK7NpuGMJY
Yb8gXqSkZtbzdh1MZ0Q8fk2EeRzGrGB76GpBz0+Xftv3niIgM4jt2MXpGfxm+q7PyHaHXxINHImT
8Tic6xpW7SAM32xugHStnIpfQg8fwNlFP1sBXTAoAMFiOm2DpKKhjYY07cRYtJp1PkmhuQ1ZGR52
HBgKwaHgWsfgjSRaX4IMNtGI873LAgdYtAZGXEGDvWRjCUzMgQLzbX6ntF7/2DQY0i+4lZ3LMBiQ
Bmg9Hg9iZoh+qzpTz49fBaTC464hT5kjbSN3k1enyNBKPpmDDS+bLwRYaKAbvzsyGAjS0T4NRQR9
z4+pzfEoMyY3z5Vb2HokTnBcEek0HQcBWtp4ezOL8HQKEokM0+HlbJ/PCqAbnD4U98V5XbDPSo1w
xWYyNeaQUKtTlTEhWKJGISHu8O42IfD/gDofu+nUiJHtDbp2/Gt70eqwUui4p7KZTYt5E9qW7/4v
+DV/3H/K8/Vjn64byZc8gfPRTQkEZWX8xT69Mos3DVrQAUdHNApXnVlJy4PnvZmYuaUOs7smLS6s
Apx3vAne4QHjIm+cKWFHBt01Whom+U7q0BN0etf387j5DQpQFADTPBZ9TuQ/xnBBNHtxAZariP8Y
eDjKaHfl6bCA8QR9W0RLzuK4OlUY38HUjjdUVUG/dwXdYjjsPVllC1gv6+BbNljJz+hvwCGUJPUr
VbBPo1AuiBIFOAeDxn6FxFnmqBfIbOJoeDGh47L5SLy8wkyeornLIqHc7+6eFt84u1i7abyrxfgy
FGuKtwOIW73vaXB1duhyYszh38axmeeUM6qfHW6cG/5QsSF4G9QCilR23yg5Z0YSfae15W+5basb
tVH/iO37wujcROBE4Qhr+XCsFHA1tSsN2TJDD/51JRBsweCfsTkNO/ebXEeLt4i3Nj1dnBJsEags
QUKiDWrZyNIJC4ZDdBGpVHe9XCCF6VSLcpJ4Y2R70wipwbqDhQzjNlkoUY/aJZv4tJcy6Y2uTwIV
uRJmu5r6MY76y3e7Jhtm+H0g1rdzKbTx5xiJ/FQkmwZyOtP8kwaqBv6c8zW4SA1DHDfrXQ+BTDcB
Tb2aMenB6mAjusz2HwoFb/Q1qqDO3W7/X3WivSe9y7gCwam4lqqScEPJlUFxOAHGCqyQaLuMH+9o
F809GU/Kq7/nXDI0oY9AjmawSqxiCBYXLeX4lxL521p05Zj/pNtAQFw/f0/s2iWITufM276yLw4m
bpWQV1HaTa0knftmsIJx5KkNEEKncFeTjxcN/3hPQfFQGJKJWPX76wsEw0FmH6xiN28KVRWkmjfc
SvjlQl0LpMVlubQL/tZaf/gpxqUPutyQWZFXx859XK1BarN+J92HcqwZwhdESweJO+lx/moYMqW6
115SenhfUTCKhVJv1VesDvAhN9Usa9KgH4HtDHq1TfZcrFE+sMuIjfU4cbG0ca1u5AYg3UqemUT9
nO8/xPbxGaFRRBJPVlKtaJQmMFddLU1OucEnNOvbT7NGZGdaP3rJnZkPi1EWhPkeNe1/TziX0nPA
EUVJ77VpEp7EPDYE/mpHxieie8XhIxHor6CeQhDvz1gb83PvAAwjgUtB5v/s2L7nYgF4/pgPExh6
vhusz06frSpx7Dy42eL99S4wsqzrcVDjH/OAe8yiTAzGAa0qAusVU3nFD1kgfjzgQHlqrxBNIRth
DagFcysAogPJZXmQKLKVHnJVBUw6U2Ykw0Tpk0vhgD45CnMSM3/jYiVgFmMDLZBOgrom9iUO4mha
0kgUfCRiEE/uEtfA1qlnsEz6QJQFcFKIe7gImmFeBcl1JCvReTOcf3PLsF/D2E3KBbD3R8UfFGp9
43y611ILF3YVP1Ao73HVE1VfA0LKnq3rxLmbH6OsKia06X5IPwaHqR21wNesFhPiTBFa1D0AhzUP
iGM7S3qjHVhIjWikAwgWyLpRI08PxKdwmUb5ImtMf8JTD8kR0aKmi61qfsFJCuKZgWPIsV2a32I8
8GreUb0Tv8RkOAHhikQUEP2PtYfIcAHBg4KMgNI/qk04x51cf45RKaPquVyJK21Dp/NNUeRJiMTT
Df+obF4DXXWuHdwv9mnfNhDwTk4fS8+SJgFfWoWSM0E9sk6U5+5bK+aUkp+mqSJawq2iSPEtYjYz
Vu2RxwQRS7oqsRkKY+oR8Trs4tZo5UN+tHLzVs8D7bn8ycAggBbE3wfOJ/kMTGQktEIsi/ajekRS
dueYYGf5ejcJKuAKE0QzcG8hNdStkdU4aECjT9oib3WDzWjoBlKKIAgdlJvHe302CngdP820t9XH
6I3Fwua+38rw8kwrkMsDsTXwALZAdy2Io5ymTAavllZu5XoOOh0+NfBEe+tM8/DXu3qHN4zNtvyP
kObsUqcOPpAH/RRZEzHsXnK4g91lMW16Hpxo77pWxZCq4UgXrFvAToZ3Qr3F3c6kqAcQctCX6YDx
iDy/fbOXH/ODW9P1YlK5EeHgyZsTzwTDb7xMv5A8fkfxMdmpWsJXtwQ+UeIWSNTVmJarIuzQgEcA
wdqj106YK48o3VCzYP4YNgvQvNz734VRvKYs+6qs4HtJTiKWenFVjpz/RYnJgRpNb9w2KmyKG/xr
BrJ5eTC+rW6U82zPwGbRSIWDS5JK45YlYntxuYEPsfYh8662O2OzvAfZvY9kCnVodWhyx23qo2S5
sNE8K3cSXOkZDeWDU2MTf2CXzhelP2HRZmnjggKYvNsdiIi+pVI3f63uVHAFk9RbB7o4KAprlRkO
d+qT9IknPad5YRTGB/e+Cqw/IBCI+Kz+rxj8NHxgvRKNBmQfYZTzyaNSC036JsOfY8vDqdxv+gni
LoVpeg+nwgzzp2g8UM+zHspC72LitWYN/dLUN/uvv5iQpTUODUMfqjZ9bf6GNzwSS3MfvsG1dMrm
a/ldxqse7oNnm0Dzrs4pAIjq/AmUZyCBNR5vZzSLAyBlwWP31tjyggUeSGg0jxxqW20qBf/5ogH1
mClEME5yMz+c4feJSbazVLzZpuGYDqeTNJCPd2HiyT9hXjLcJr9YeNUY73a7lojRrqoS7IgLD5v+
JyepTrwZ5UXOjWGONZfJVeh888xTWOYAj0mqKMI3m+fO/xxBkLB8H9+lkEH1OJ72ukq15V69J0Kk
mdck3v15KXj79HyyLSDsxctJr1aOPYLJTp3ZseSBGUyBvKOkCWPgqjrQUJD+gaEhMrIWWZt1z0qD
nfIyGtPyeCVVazAEDAU3XDYup7uNA5HLqI8Qu/+uMUqeiN5sPurVgqzgsR5Tl0zYBfuVdBQetYT9
vmD10/gTliFvM7uDZPDmQxTXpUMt0hp3LLkCiM3omKYMqgpOKe10g/lNJq8OeRIPYTKaf3Tyv9R+
ZHJwVne2Q7pGVOR3XnqOHZS5VbVaUxRBxwnQDqGhYD+AhVOeiOGsnpuIdrPCGjsok78idW2iI243
lVmCGB2ekXnA41oUe5yN9d2lXevDVrfZpC2ZdGIwxyQSBAapl2SDmAQ7sN00hf0FMaumQYE/u071
zXOipbLEQa6muw7pbPyMRO12q03qrywGtQpn+ISSYZAQdKmxMOgqEIBViatI+kLb9es7bW8i2PLW
72nOAbyp0EfUV5+XAXpO7efUU8LRY+yAH9jvFrSaL1XbBW84F3Ww+BJh5n0BEisEygJZ4oia4j+u
KjgNrYm608T9W/55U3reYC5eNfTdDE3oH94MMS9fr5BHY3C8lBdBSW1/CCI19kwz8cGiliazwxnb
loxDq/dXd0Z/89dfbbHMH1iw2/3uBlNWvo+2IgCnNCYwfS9z3rdMpnLbTs8J3PV84aG9bVhVJ/kd
V1+ecVuPuHoXznOt04ypAvSkf5Oazi8hB3QZPndXp6Erw+26m6OboGB1M0ns62RBBEylw4uHV2wv
h/EThGwa2Kh6aEC0O6JKRBJs1ABPlWutwXLXUoZdxSzBsho3snHTxLKON/bIXP87ghhYtiOeBXCf
W1HVStrik8d6pO2knpGwNeZQn5IvgKFxYBKmMYd8DTqeqG3e23vHZKyNq+VXr5/xksyOJ2pDOA4w
xzk2+FVbHTsPMVMi0qy+Wiike2/nBUMH0dKaqz0ICAV5QvrZX9VtNj0fCUCg+yK/36xFcFIQ5KQ3
/BLDyDXX5hMrMa5Z/OBygg8HslP9TYjzvejGGANkyMMMUMJSvar/J5HBlksyEefAEV4BtKlJTGXI
cFzfDo+CnwUilCI/Ffup4K67Yt8DDs7ShN/o4iabUhdsWZ5UFUad773tvtpt92XOHt9PdEiLq7PH
PvNWpCF9e/KIHXU9C4T/1YE9HKSkjSQgnRFowcnNmnDQQ3Dq76RcR124mQ2NLq/49L6WbHGCI9+V
acMMXokQUmX01Lau6KY34JtGGkgx7DrqHhl/bplzuyXZ+7alv3fPQse/KrA0olC6DzN3Fgp590UP
wyR8Os0ppOXqnpJUQ6am/AYbR9wQta23wYZk1Qb7McHIyyMbi6cXJLAUFKK/xkOPgKiS1mqPMgS2
D/l3ww7awXQNWLjb8GwYhmAmClTq0/43MxPXg8bW39K1erT6SzTyyCU4NGo4X4QdLkCRKsFY2iMq
KfkR1UUKpQGBddfPIoJNQ7yWVkQ+AATHWOrW4tZ17mq0/xFEOERoIlUNu3pGR3xsngh74eHIorx8
4tUsZ/tL/IxyFzuGz6kQnwqpRji9A7TQ5kRiP/KlGIyiJmdl4+Ebtfqlq8xD4Rq/X2yuxXfYNJeP
B8T5HC8mvTryCQBN5SKTiLNuTX9jd1NZ92Tpv8xe3cl+FdpfsE1Ovb+f8D5M7CTpWVGHFoSbpWmT
LWpMaXbLMcXKAW+Fpa8hZ7uopSM6WXFKJpLyqAPgFywRcY3WsK/3pIeCMfPdyoOezrTXSV6Q/4sH
/xeiIrxzFh/me9kF1ICnGAnq/RPxLE3iUEnLk4t7l6JrlF3Tke77+GlFZ73zMmPgcySQcaZEHfk1
UGCnVUZ/nvGXUYcw552/Xsm4L2r2VLJVaLwp9R8DjmaRGXG/XmUh8Exrl5PzjqIKqfWy60e4subc
WJIVakxxrk0pPd3wyDSPhI8P/yfiBPO71iGJ3nf8tQiHdcMLFVLcBxL+aRoLSlg8hI9Vcj4xPtKv
gzhbUaEMNMLPjY8OAm6SquJ4PRIoIgsGjw37561fHfJHEqO3gC8VweizEPp3goYMLnSd0/yLNZeu
UfkJRGKInKUov8rUhGRbGtLqUzSRy1nXeDfpF+dcEaW5J8a0JLmL/aDQ/ONYuqOWR+3c6lBZaR3M
s5iYn1eYlh7bSaIpKjrZSv1oy3XEGABcJ7UNCX/1s7tGIhtAt024bRl5IXQyg0xJ/tL1QDzc9PwH
jmjtJof8R8HCCDFP/c5A9ZMYr2JkXxfvH6KrakrxxlWl7Tc1jDi/P98QzswkzsYLYhLOan8fRdnp
GW4Fe3NjzvCMfA80VRW0kfzta5wsP3hU1MjJQBYEPyUTr6tWWABpJmoW6SILam59qngzL8bbXSqR
t0XTlewHUcBg532NXBdqwGsGqgGvy41B0g54zsmwCTsLd0Q3F58NZKKwEDC573MRb13Fo5ncQGz8
MIcizIHsk+XXZVKVeOdUnPU2wVxV0at7WjorSqPBBYAKaCDE5mStF4IuUzDhcFJLe0OoOc2w/xRG
kLLLt4m0v2j5XEhldNDSvS2pAmEe0+iJoCVcWxWpvd3DX+RPWPZ1OMMV9asTgyeAOPVn0Kd4TnTj
51gqSvJ9rGyLaanV3SoHPr70dCG8fjWR9Mzq7jJH0qOhNydQziyVCkK0wHXILK4LDeRyOdIR7i/1
L2LOdCOudLOb/cTg97BCpkhH4TiVNlpvJS1IBniha9NHohMopLlmfanuCxGlyGlYjGtR78PqC48v
6C3wDi6DzugaAbiAhMjJafU91Pbevfbrt7gd+6GCCVxa6q3jWBz5jqNLdv1i4w9TR/RYFe+jIvFe
esX/4WvZj4swAX519lt8rw4mxeZgBPsOpGfFrKpm41HmtbSEwHnEAFw8DcHJi3tH31oAlp0ECzWO
brPsQbsHUrTY5VQLQRc29UV44GRyXsseQtyfwBHLqmgcOwYhqvSJrFTZG+ItdtsW6iAENjD1Clu0
Cb5oiR5/B619E3mr385oYkF0ekE9Rl7rLH3M28tHPmRjEoA3joJ0OcFg1dKMFKAlCDMbvMKK7N15
EHKoQShbfK3SUjWJrxXduQrcjjfb70JSR2iXzP0eWsfBlCM2rWqRxWL8nXzQvKSleVPK2MNMPGlr
Yod8QQnBPccxjcK7fiVoSN38RNhoOAw0Wo1yQSxbYvkhsg96KjGyOwS6qWpLgfhdmKcwCmJ6D/8G
g1JeSzF/TAJM+VDaeF7q2awrStPzNU+LAVrGNRplKqrJZt/Y1CcuQ3TA+6t5zJAyjeUsHOOxKDIM
RO6zdO2+rsP6QsBt929TNI6UCmyM/OdgE/AhfrSmQLwZ5KTgdRLcW0MeEnUlFxPfNPSJoQW067+U
81zMrLFlwhWaNG1yGl60Xh0Pv7GBKvseas0Kgs7BRGtvg6eG9sctEMJyU0SkHnasUd94qk7ZJavY
/x29+zA7gnYVPVRbnkp7jGQp1NfwWF6Uxicg8c2D/zu285yfulYQvTT1GrGg20/YHoskYOCOgHwe
ECGkBUxx/sodc90HlsJ56pnP7YLizqjfKtoPsryVXC6vgGr7U9/l2rasG+4OwbSiBVkURthG6W2+
n6fdKZ6djOqZrlfQ/fgSTTDcj58jc29mEnnDX7EouLqJPG7JKLjqeJO7ir40Id1Ys48TIw7T64uH
cAn/E0e8uKMA8TE5ZNtp+dbD/+kahBK6LZD10Ak6CszTMujE1NhhULQ7EPb5vlqVsqin4Q/IyCI5
OuwBKIPLpy8i+a2eBRpMZYhJShzWeI3abo1VqfQoLtZibS7wsv00zeHEm3u7rLhfQnLK165cb7Af
mzD4KEsphUWV7RpradELhTe3jJJscCd9Ko0EgjqglMktK+z/2qKDOsf08o8rhv44BVGYJuElXS6m
G+7uETjoKFtzBc1BPMSGVJUeZEEKLvLic9GK/tBV7QCmmvV6V5izYUbmjenJxwoZJbBGq0jw+our
roRnlE8QQtT8hd9yy1ksB8XsQI+qdK8v02iqSFMsATrH4u2d1TbS/clSomPajiK/+s/2im26tx0q
jS1jIQaQOrt0B7vP6X1TalRLte8B1tkH84z3/2QHBagB2SZLT9KiO6dMeLP04qAnyV00zw9uFnaO
91N5Xzt7OChuZqgiYYOqPsO4GnaYroHePXk+IkrZ/3W87swtwH9V+r7WipfbYI+IvUNr53yfXZOH
f7Nl/hStEryZJof6NwYRGdkJ9sBv91fzVFSMESC3dH0SK4oNWPCNA8vM65EW9sbOz7LKBu8vpRTd
0tuU18dM0Ezn20/Bv/5+MAfQ29+R92yCqSCaPWRW23B4OkVyxgOPJuF2dQhpe5talEqg4UiWHZgq
l1tckuyeE5NVz5vKNZYAusWO9FMVjdNh3mNRXtXK6sEgkQSmKaJ7wi6/j5/xWSzdFOSAxw2MAvUv
VgmoF0ZOF+0XxTs2xlFdmEnwYDm4nUsw3xaXt+PNp//T6ifxMdwM6TajlwidA2TpW+q8RlgpCGdd
TKSXpPQy9hqWBQga3PC1w+EhCbhwls718izaSDOK9nU39OEYiC1P6NKGQnPM9fW4PJOqgAJoN1P9
n8XiQ6D/32dcnQC2R5lHayxq3bqsW8Wdc55P4Ikb7o+ldbtq6a4uLt6PQL0SCBXxXW9v9nqcKQ9z
TCiPWDbc6L52Rj3mtZkP4TJ2nsaXRpMzGp0Dnr2uyysIMkx5AZa1Zb93epGOLQRefuL1dtEANdYz
ycamQ4FDMgw9fbEdF3OBo+eL6no2KGOEOrHKvsxsTMG6MlhoWqA4RT6fmDapXrYy2Jv/wCXqiZzP
cpqkO6BgDrhCl4PcOPwQO1GRf2D9ZZaXjS8SFEWvTP3DPt74aeIKVXALtAOFzKVIWC7Jyl7JC7eK
pfo1qTgRJpkxniausv9cDQuer8+HPFE0UV7Bji507/6VCeC1n7Fg3crv63FeEI0xJWLTqB53+/V/
CVkbqdCRJbi4AYumcJU4xBGLMj0V/t097cfYB9cC+qI1h6cz0ilILiOxm0oXskJci+dDrPEsEN4H
3hAxmWhQHCRoUR1eWF2QCG5pC0oaSQgwsvctsWI7bu8QwP5vCrT/Khe+7inlP00xr0DudroqgjKE
fBeIsN6sJY0c4aypWRjBVGIEc2quD9eFCr6f8ZDC+eouq04Wf/frUvPqRoBR9YVcChlGVA6dW1mp
XCpPNJYbPXEykprc66WdrG2aLH4x9ljYFyC+ofHjSzQDyP1rQZhSu5DwYu0qwg84+OpDjcSVbyYI
4kovHotBmcap8Fr0Yiw1IyCZXAINsNYTXMrxb5JXjhDozK2yi21KFbfwmOsLCFD9Fyx7aGnDPI11
Qagnk71eNtBMzzCejM1xIAbP2p6KxgPeq2H5Df4RL3NkFLaFPzvthHqUG9oU5KYED9eyPpks9WB0
9ZVuy9ezOgmz0t1DkH4iDBaH8bcGpDb22tT5X3oSKwFR1XAv9fKfgdts5ciOJZBaTHHQCFvEFLjS
vxggi+Xwr5dpXTCls0fWenG3W233JS7G3mDz4Z+p5Kp6xjDo+YUD36ElNFIxETxOHItX/R4elEPD
XbQRyX9HcC26u2aJluMjzjOnkYGY6Tl0VE1q4Qa45ePf57rVisa5Nq2jtiTQFLYjgp5lLp3Hzv5Z
6Y7XHyQJYoC3c0tlqjOao9CgTF8eCdpFQiUppx32eiziwd8QSX26XyqyUTTcGBDyMP/SlZB9kpQl
200Kk34jYP1qZ+CxoPvXhA+pWQ/9X5pZwofbN5x2KDsJDsQy+5Rfu3pGLDvwF1o/Mzrgh+W/QgGE
7wgu6qJm7hc3E1M7mokfMJEIt22jUTZ+qcc1a0OUz9RL+Fr3sfiM2klOlLgmAQtsiuhjCSoQlyOD
n6UXHSHxa/QdaCdKrOs+o5WeRv0rUnHzdaEYpMDluLJbIOfcE7sFl2t9GOH53RIywVTN+mXjVKrI
NuFa3frdDtQdc+XKc5Hs8QnYMHO5pmYqaWW+s14SLJ13jYXQ1Itysm+Vr0ohnVndjqSA5qpdbNa7
zjw7jjZEovrmdUowF0/MLK6ifHMZdULO2BpzKqDFzuur5jW6yw/wqfCLre/nOMRi0E4t4yd7TuGj
XpIW4rYvuqioUmmFfYqb+41eAdx6Mih/Px0ru512+5cgfhVBGI1SqUhuuLIj8oJongOluzEv8FIR
zK+Sj05HL55eeVsEi5EGEvpBsav+kHFPAhUPqrNCHaM2/6bPH1QkWKrhW6QJSBlPgizwUr1Fmedj
kqGtq1iEguF0NIAbdWOvJOpeOSMNH8QFAFZgL/lwk/XBSDSccndHByNjEaRV36pY0J/I0XdmRFEv
LVJ5IoKvHjTSf0s0dOKnrA9S+PncK+KlbPG/4NXI8Ypepn6Wb5+zuuojpfNn0GEibZMBmq7LMwKz
Kt29cTzX99FxQ7CAn/u5x6Nk7vadTFRSTgwlvD6z4/1KA2xMy7y4Z3x/APDyYwol0zTraHsz89I/
LHr0oWy+jAZsGvQvPMXCcNsdVZF7uPSGVDICK4EcFIw3ZjT2Kks4jKDIVO6JYmt4PqUmeK0Mk7nw
+NBUElJ6A0uKCPu8gTyzSHst9CWFWLeG9BSqLOrONIaXMg84u5hpkYB10wUwnlfxHwWzW2TKoqQw
K+xyJ8ymrxI69QxvFoztCfgO55vDxEXzFa0AruyE8jDTDzQ+IbZ1/57O7IlmJ/t5VbXFIisI2ZHk
oo9tT3cVuq6bUuN7Eq02WRMUy4MklL1Te0H14FHGsx4A+SfoXPOYFUS10n1ruKukvp+hauzuMGHX
f4wQfajJZOqLsfFqcoSz1tjmm40zvyBIXlomjP7Z45fG6R4+v9R4Manyf6rCEZZndVbKGD6/yTMf
rbEqmRn7TkhGGq02CDrW6gp5ck0MPjyjUFlfbH2DavZDYylfMLs6Hzk/PK/7sgf1w0+i6LxiKvFp
3L4OnCdP2RPXsxwNkT1kVgyRYm9/Q+jbvQtQ+oYqXAxqSNNx30pPjaaCXIfM49jCaxgJpBNQjIOX
wtpWujJb6glGqEyKnxwSidjekmyc73EXsR3hjF0ITYI6fouNFR030UQneMsXk2wCU1RKrbTEIc6z
di/O0k00t6DOX7xvoVGlMZAmQLLb/e8/x8iDbTP7LTKYEXA/JF+xfBzto33w/iFXI/DXGV0fRkUC
/pyH9EwbWoM8ndqfacxe5fCmCv25UnOLixjYqyVR+e2VAF/1BW16u7I6dZK2dN+keIruSMtq3VGi
93foD6ju3QmM66Q+uH+2zcEl+FR8mDGHwAKqKSfbAR8o/ouwtzVOFb8TwzuWSdP3U84UPIzFywk8
H/z/Ki2Lw43/NcO0SJp7XRRhMZPjacVLe3059hgRIlbRt7ttYDYxAuQYb5+p53FQGFIbooI02ODX
+22QSV7Kog3PTJYqDlTDOFuoB6kCYV5xd4josckgX+L0xv4fIBvhyxhIgSlH43er0Bu74lBaEC2M
dFDVdJU33aDQ4cN9TdIs+VvV0bQAeGJ/+Ohcfl1qh1HWBH2aH1AOEwEHS2tPJDNZT7obsz1SNZzX
9TLa3g3S3QSEPtmVhTyFp7NRj+DcTKIBsQYVKZD1zfmz67LU/li74jucEcD/xkyfpyiv2ecEBNmz
75N4M/EEnMZ68acx2sgRJewZ4OjMlD4ppSxlvl2cvr6cnA2ZcAuA1KyqKtQZq/jntVeDkUmamCvm
XBHXg9AwaSLN5uPDCJ+BfUkiyCEEEB5cUhScdoBpjTFBG01F0Mz27ZkAgDmHR7Tge5gC8NYt+Vzw
31tXuNzfDpQdYAExC2qXZ01ho3hvqxfYB++z9sS+XhN0t4595nvQQ4obmZvOwzcEKTy9SLR2CPxz
LkhmpfYAkN5VE+qlXf0+nWmteYldhWUT8bBuuTScim3ACLtOjD42hvzJaLsc5cPCYEyggOFMSLgs
oVtzw5ET5X/9ndZ0MWnQV3KbXA4LkPJbvsvbZWuZhrxkLk6nus1ZNXkdU4DZb87lOA0sfKTYchm0
3Vjllhnm+ZBQgwBd8pwm4fXStUqOGAee++qfh6NWZRvBXh4h/G+Oa8V5yII1dIEgZMNWifR+2nhJ
ECJGcwJZnwrei9TRqg7wAXzfnvoLPzbQ0oz51CsqnyagclvJK8ouU77O+7s+GSVC5ax0BVQbr1Xi
zyX+GHgZU0diyeS55lz/dfpLUcp8SfOh3b8QuUX7nQiomlkmCj2bY0w0/6WpyREjHiKdswIsiu6z
/Tozy3FgvxCizawfck/gkY1MvCKE3zhGDH5H2sb4bf5esywzn0XrDJaz9lekvGo8KEdlMQyNUEMz
czV62IsTYcLl6EwBbf3MXQ2ha/jZUWX2VvcTmZPWyK54HHEpoO4/L3xz/T4Uh5wvb2+ci/z2MeF+
14pmAza/d2xTAxis2GlcoUS07TNvV5ly30WkC449Pt70xjivhUmFfy9EOymQxKxUs02ntJoSC4RD
PTzhTM4dg7xgDFQQabz0e7Eab5iQuV4Os3b0NbGMr8LDngx6MDtbDaxsTSHj4KFuqwXQdO4zsw50
aB9uKvf7TqgMUiSiR6QZXTZGHZEJw0cofeEMGuSEMeDqsB6zlgm7KHULW7l+PDSMFRJgo4LBpCt8
Ci4ntbASRc1Rqr5GOOaiY2W4g36djN2Wlgv2AWhZ7LdC2OwV4+4qPWTIa+vDECMOhdE27Jh09z++
QVeDHt+pQKl1/u6FyTSub5+BI+KUGliS6VfBrQmEyefxyrW7wV8gI3SS+1yxUqJ64Z4jK5XPNSrn
kgR+jMWs/hrdLVDpGOP93Ib+rdIPdyoMGOsSlJ0bOWELERnGq8j3/zEt7adMT9AHQBRiwkN6xhx5
hjeAAHGIcAqgkPvO5n/0iV//MO56t4SFL6QAwZkj8iUrrJIyux1IOnU1hXA/48nPMV7e0QbIFcJA
/sHxiJEQC6KI/mp+hl+KcZLtX93oFIafg+sBPyECMjd0h+y4usM+6Guh3PafZ921gS4lcO1wY1mo
ni+ssT0JaEiMxX6PUApWjl4tP/ZxDztUeWxxfw2T0cBhN9ADVJmcRj1UP5Z8ON7X56bGKwD8ooZF
Lz2Ai5hOeMHGADjGYEed89Lx1mWgDhUsUTzF8djtPVbPYvpz64PMxVL45dVnpNnD7bunN6eYTZtW
urFUNQ8V9JmYqtTn0TNkTMj+/si3jjQOUB/UIt1UAew6eUG8U4SzYrV1LMqKgE4qao353RxjLgcA
0virykMd6E3KZ4phl4K07UOm/eS1ZBmPuryRopE/uZTSdBYR3QGt/Mz4XLeGUbJSg0IAOv9drTtf
Nv8zPwx69COe6e4v8PpBJw4k90DeTo1BiIYPNAR17hVTUfXmiC6tjTpmvHtoVutr31BHhL+CTdeo
ymxLfpU77s/wlobmGkNgtTB7UdSIBkUyt6JWrBMhVZjdyOun3xVr883YXRzPluk7Qew58f5IvtiN
y/bM2DO52hV/vzb6S9iC8nr8PNJ25OS8bqoBrc7zlcpxQR8VxL+csfdELUSGicG3xKHxw+8e+JO8
OeIrFBtYvO5SdMquvstTBnhsuf9gvCPKcUawW9hKrMPJGo7fp88LK+ZpQqsNgFSRTIya77gdDAs+
KG9VF3raPTYTPmdIKdHv5AD+0sZmoGMPFzVu1R/QHysmxXVy3OQ34Nb12AHmqOi9L7UzDPqRYi54
jYbiN3f8z3KODzlNozRyvEiIdmHGZtTcdqtXEPyHLNQOtE5HAIcKw+anAGi1UT+Ufd6dLae/lPR7
YAlRB9FOB19sSsz2/fg4CmqVMoJb80wPN6krhowEWP0jxUmW+hm2t4dFBT1t9jRbIA4SXDeJ2bg8
pi4mPyZFo4eFAn/GPwW/nHPnjRIRjM+sqjzVVN82MDYkn9tXjWUrsMWvY8cHVJMjOdkaIRD9sKqY
SoDdU0c8OYL0GOq+BSQzfjldcx9D93cs8lzpC/FuEwXDf5cf+5Bpu6C5THx9sbRxvq9jMMs1m1nm
YyodsvOvDijM90eLIkYYnUXWC3/Wo1YWfJgkg6Us29sqHMK44Ad6GrQSQ/0MSD0cRqord4x9nZCE
WGzhNCTEbiEQA0V/iQuotnjetaHKFWRruzOEzyjl9OCcAgNnfbmGEd79zMYO4NUsu8H4/lfwnYy/
hUuGi9OuN/iH8U0osY0cEsKeV/w6HDo5CuK+u3kh17CR5OlcRbtRKF6ZyNuzp+gTum2AM9FwWUp/
oYI5jGix7DCKiLmx0c0d41T+ulJ3fZTQL4mCSmyR+mu/QoCThfrl/rBO4If6pgttbxSNWyhBW9Cq
m5bNnnoNS/pvJWmJk1Odimy76Gvis3ihmvhhx8YODLFuavkBRdnJTpiwl8WweH2ipZs6GAcgepcn
Ph1BHUL3y3t2Cg6ZwfIHtpNCMtVfOg7n9ZUc9unAL3QktgMcY3/ExopZvRe21Au1qaqEgOh821Mz
OE/GXdcqk1V+cQFqPlPieo1WwRYL5XgFrg441ljiklIcixgus5D0fe2b7TDLR2vCCb9Lzx3jD0NW
ZXBxxqBwnloUBrb/N60zd3t4fN2BjruUpVvLbDS3RMYq/U9bglX/KOXL7aiU4thAdQfz/UiC/TXQ
xLzSuC3mPSZQPtXxI+ypCHP9ZyXZIT5fifRbNFhpFR9fFTrRaihdUyBub8Ove14Gjg1v+pwos/TF
FElsceiw7LdBVVvckoQEjyEGL4HJyPr474ydyVcF5zf3jRgu7ReX/Cu9yndsd4zropWq8OXse96o
HKHk3/GmdxIx88wfS/kowKnrya3USh6XG2Zt1Sy0Va7xHFGWDPGOxTg1HwzntFv7NignaS1rZABe
QZaInZ8QsOR1Yy0mxKNsk42qh7WwpqJljbio19337Zq+1Nmz3f9Kg/VhZ2ecxqYMvLPKAbs6XViy
zucDZLjDRYbPz/1TpjWQZo5tpNbgOVbb+AWragcfjw3XdFAyD62A2Lff5ogI1l3cf6yNeDh/4bzn
HrYaXI0X5MyD5sRwv9wLyzB7A+Of2hmai9/gohKvk3sw8cXn/5Tm2mKTH7XQTeroAmxfLI4/Ww0I
IphulcRTU+MIb5rYW8i+gcm5MzVIroquxyhPa8EpcprT7JPSP9RWR8IO2xVHkydUVKwqmrctioYm
k2Zjz+s8g33wFElUJ6f2EaCUFJwc/vraaKdFSSspnjjqSY8PZCeuEMpLsPDK0Rx4aIQHM/8fQ3OD
sIb1V1sUl4rmfsM9KNb4aKFJ0SfWK7HtNWHxPMrw8jai7jYoPsa6EqpC+/N0rmgaOec8BjuiUt9G
teh7zPjCJFmj8sh30uz+ubscoWDW0LVZWigbqqZL0PucY9vwpg9H5EOu846JOSpcxmD+nSgCkmwx
A5OfYPtSR10QecpUgf8PsEZlU5CV8KT0Z/JEa6ZCw+EkvUO36r9TuT3yScNRrS+uQKb7bYHn/Zhn
+nggWpKzqjHjWSxT7OV/VXQaRAvpu2oaK39oogb/h68C1Uw5MT6rta6ZTlhO1Gw0+2YTtvSigSQn
oCb0xNcZwGGJK7DUY80UovKSnPHbSlxJL7x40thqTKlF4SoQ60JoNWRImukaFUBv1rAw27s7G7M0
SOmZJnBLdBKhrkBkOhOspPmmQijekjDIsC1r9I630HYKjg+SxTxl2kd5ItaZkypX4G4Vmuiw7Pf8
hhM0u5LyUlDQ/YuCxtDsRDF3Rvfy76T/x1qYLzY2XBBoQ86q5/2XD/fGnXvyxiGU2vw9HZZJF50a
YSZDKPHTiyqXOHSp1ZnM9eZPYU+h2/oSfy3GfRiOCgmufh1UdWyI+SiWTZmhhSlyB1oqwZQ+WiUQ
wC7/Fd7yzLOzmvPjX25aE2WjoVWOaek68NRwHvzDR6pRbxoCi0F5z32+r81vhekLfssuYNPrXNx1
Awc/hQRrQFDw4wRF8QwHlCeDwcD0fNjchmemBSZe5xC6943rvOtVBrWMIG6XyqkyPxn4l0baXufo
gMtrBGre9YXIaH02IZtfrNJ3Yq3CtAuPaywURzzROWzjQ3Rpp5StFwlCpzmxcZAP4OkBfORmea2T
7c71MhsHHcqnR0f7Ovqi75AIosMSYH+ULwYipAJMQkh8HkVhTGn7t2DC16AOLKwAMbXbx+Yy4Dyi
kn+KlLajsJEJpwhcI9785OJ6FN7Cl7N18C8QWIU0emmSNdM8pyHSTPwYilforzOd8ZRDKag/UCz1
jRhu2qHRb0ct7E45PayWSNAxAEPTs27oicJMf0zXbK4Lj9Lo8AtecJo7+vrQ+/CehLIYgqEQt7jN
qxxv6MyJVDBS9gv0Vh5EGStksichm3SbzSAfERFJiPohiF8elrrDeEWpRedAQvSlSR0yfEfjy/w9
GqLLbIL0nhrXend/MEgMnbGA5+TgqBJR9N9MeoGjzKyy8Ip4g29xgKfS0t++j8TEUf8qNchy9yJK
sTOmlhEm/5TqpspTqiPvDIb8zfBXB/649sZHLshl6ZB5Ibti9Iok2AoaHzuP1yT3P1YWtH3LjTey
wuVN2ZHS1iU8EHIjseHUrcO3vqFSZTUR3ivzyADluxa6RZuB2k8eUsdTYGnenWqD6BgQb6llmY4L
gWLITU+zhtxoXhamIZmOHGsO4YQ61S+cwIyJmAoEzBG1zDBJQ6nV5OIhkK7AEwFrlYol4V9XNAaC
2ubv4F+QP+QQOEWw/+gc0Phh+f6ItcSeN9Uy4XblmCH/lOb+HAOIDwqI34Lxa2WSHIKbN9tQoCJO
QiygON8dCMCGXOMt2Bxkx1TNrRPTNjAGrGgO2l/1i+Byao1HoeBcMzIlyjU0TYvUdJ1VNvfgTRT7
H9KWWeKJuPWhFemogyoqLnxK66RgWo3NZ/TvMtKSqDgXBB9/LH4rGOFVYL0CmCNS5IKa0UptXqKH
Rv02KvCNcvpcYFGBwFvg+FNzcTB2uKQt8uz3/yJGefpm8PNSaRvloc6o4B1Dl1XGxiyKeuvnWMjl
VrsFy2mqARMLf/LoCQ3benP89Z3UNOkuZIND5wCDSFQN2MIyuz83iPqX5zFaW79Yugn2zq7hr2fo
KGifjUF+IN7Dlt1998jb2uP3M36oJRNPR3heaFF6pbOmKLuYC0C2wFRst+n/EefQBkn0JokbAui6
H+Kxd+YDDmu5GD/5hNwTcYo75B0d2D7dQ2mUiAoCBjqo3BlOb8N75lV/8eQykrrB4CsJk0sDpSdn
46vDESdNPCk39k1N1yYT7Jw5vhyP0ahlWtG38ZxDs5DXFQpUlmESx3SCO5T3zej2OCRqEieVotEN
9mN5CdDW4V0LaHs8JEbG9pnwUmt35XYVKyL1+fhz3xeVHGhufEtRHd9+ttiBemNrodBeOg02hGMM
6KMpONfb+ja7uH8YNY2cHXEGqtMSzv58HogGAkl1/EbEwwQ+fSIATvpjzpyA+ZEoVYIJGiao5bhB
AMGWxSOpc2Aeh92m69k2I50OQwy/A4h2iIsOCx5Uls6/Q872Jw4ipzlecZKZ6xCa3C+46XoR7L2O
p3OVgEv86hJy4Ze1XFK//mk0d+P3P2vsMha2KQDPyGXMpOsFOx8qkrIM6kQ9WWEwWqtKJUePy6lP
Ls7wdY/js+Mi1EV1qm+7A67lZfreFzOduVBBIGaY73ZhXsYM0jn4xS93pUGFzFxWGEtcgcXW8ugv
uroQOZi2UDLgsv7s32YEBtdWtqATBJCxBAuP20xDqmm3e4PCiR1T0x0t04LhSJkW/J8BY9moaUbl
ifiueyi0TmieT4rHu+AEUX0ullxNZcy7Tal8TAkZVmfHfy5PJRwd6FmvgZdX+r74TaA7Ox+HH3+H
Hab3cLj6YaiPPzqXjhVHxYFxa0fZD3cNV++I3Hy1ny6motk2eGla/kF1yWgMvct+e7+sa2oXOreD
r6ZFZsuQp8PNfH4Ithr0ZWNdU0r0euiEzgyC+r1548SWnK16G0N/LFDZ+sC6u5SOxm12bM3pZ1oq
AxwxTverdmILYSRzRk4cq9ilutqBBDXEqnp2vrQp1Y7h0/ag9yLCaucH/RKTyAOGjHAQnOMPAxin
i7+GprrNJlfdz0Iv2LG5XSQ9JTxWp6XarydLGgHLvB3TjzMTSailKXAQfpFwnGBh25U+3PxBirnA
5BovMHWhYq+64byk3wJ/WCqvER3msd+fDtozIwJMe6evQdMnC+NVQllX6iaFDrR918varNCsg3OM
+9cN5pGyRvlYI1aEfMtLc/4ICb9CwAApEuIoGZN7tCoclHZ1fYPYIqMqMXUIUMgokudHTKxWmhQR
kUgo04Of4myteke4zuSuPNjvAHLhkWFmbYSB5WlVUMlEE0U2F1i/1QwoYkQnXedS9f8jbbxR40fy
max13zAnlSAa9XquuF94iIsPqP+4g17rPX6dQZZwmgqzHOMLY/Gnqsp9gKjOt8NX9kjsbmQrWD2E
5Ea/9cTonF09SVruskHvB0B0NizHe6W078ttC/TrvmY/aWqzV+IgD19LLKqqEQQBHeshRiuppn/o
39XGkzXVRsSESeWXuO7U2RzaRprchq5mN8Syl247ZXOkPDknHWcngZeBFOMbpxWF1CmAmnmWSFdk
U1M/KEMtp14jKfu22V8ULPdItELFl4qnSpn71ncO2eman88xC9Aoo3r6OXHUQx9LLuCNE9e7VLcA
3U/boAXQUEgKpwXaDvvCnW6BAgp4csnBhNWkL8bAkC3Yst1783jVLuH4yTW4xsuEwrxFLOaJrSXl
LSQjVnJTP7HI7N/TlEp90RDdrtpY1ymY6WYFBEnO9+RpVSdlGZNYP5EyBF0w0gC8VstLKrnNT7sk
SruuEYE3Guw8nz2TAUukwyvp24UhruDXBUH6bl+/W4Ho4LMTMhEnbTRFkqq5j/s6cu4nGaUzcVRY
EbNADC4HpygIiiGdCbhQx2AlX6iI6JkLWHYIAuoNNa464C8ww5aI6XiSilBokq6gbboq2u7b/ERx
4OoAujGylxDjrf+Wxj3kUngjthBp4jJ2yTEDwWW1LHLvSzQqAuN/iR4iFqZwL6fzi33OVDz9iXBd
DQFzMA38i3mGloRJ1v5BIMOZz08xoFQP8Ae/wzujBebSQvg4HGISe/IZP82+WEZ4ylnoOIESbCct
FVrbPYXIHSMOL+pHMBU8r4ZD253vNlFRdFAKs2BWyS3AagqcK/yJ7JQWqYwa6oOIh0jw0Y52WlYY
JCk4Sp9nIZBQt/yYAoYFeBUq/iB8U8PwHaWti0mGtBMTkqELfBn+zz1CQwVNBH+49iuvU4KUt5AK
32AEBEbutmapBLHBcvq/b33zoH1RBUII3utao5Ti2JH6XF8S3GCM+DGKsUv5CK/WV2XVpcqe2dUE
kSjA2FkFZ2dxzQHF/xC2CLcNBr685DgZ4Wzxw2XrpOz3g9v6safUp/qnHgBu3xucu2w8gknMbgFG
3t5etagaX1ukRtRLblgjzvHe/pbxGO55pf3UzReP8joKl843QZTlnLRN+TSOZuAm1DHji2OjZxG5
9kCdW/1HU5l+gvbrtu/qgWQAZhrUBBUalnT0p7/JAZc/OkU0fmqESQY9Y5St/OvbcJ/QO/dFe8bV
Dt2frQCGtWWn51PrDWaZpQNsw4c1YzoK2jN+abssb33sllJCn4FzE1Wz06VUVqFaCdfGQNQ1fEpV
ya2BRLMKgef6QtPhF30Hnlk3lpYxzkYrAKGTTxy/y6Ja+B1/DCJ2tRSkxsPYJAMRTAZtPg/iefVy
RoV7jub/whF4lgaI9Y6dyjlOHeFj3IvXdZf+Glu069l0qMtHLSv28Q8c1X46XxvCYr5l0UCFs3kk
dOMzRPAROA0bsBRf2OrDVuoAB5ovRf4JEZlKRpLfO+y9EsRvEX5JC5HQd8FHuy8klg+Fbl1TZPxJ
wJX/0Y+hxUHPWd/l674EA5buEnwk9ajuKVhKlcFRW447lwehIIrjWCpwqX5KyB9J4iY1whONIadr
PFUybCZvtGQCxtTpAFH2mGl5iduXC13YQndtWAZytUg9ZLoMe4Ttv9YkO8/8MRYPIvs9lUSV98Fm
NlVk+tYDlLy/5fya9VT1SM8nXN13v1J5HlGiXD5Vd3VdGEciPntrCYy4tGYJVHpQ96HDT7qtkdWE
bMYtXf2vpHHofZ/j7rMX4uFOHCsuV6GCWwc0qko8mTeVxy1HEx6fnW1UK3CESvmIfeY/STETIZxl
uA3jW4cNgZt2llssn0W97MyFTyjxDwaG57DlsX1BpyZB2dvAvOT36pZ0Z8PurGQUv+kF6uTxSP6R
RN149MQY06c30SdHUUG+lp1vJ4wO6BtfALJCMk3C2d6xuL8Dpddu4JDdu9YTkvgIeJSsBVl3J2Kz
mWjv0pGS6Q3R8lwVNyvFaz8zZRN6Kq5HhqW2+VjX7Q4SMFvYcWu/0E99vaXuTltiTDoeCWSd9H3e
gI9YBRiiWsqLwrlpuFPG8cEUTFMl3/z3/Y+0EZBztzX4KUwhOBBic5jU5TQDw2//Tns52NGZWE3a
8+H8XfmaDcEl9qIKh6zHslfqBZmKfXHnH2eUGrJlxqfiM9sLLwsve4yTZLFP+LR4ohiESlFbeDP1
R6wOt8fxW4IrhGgncycF7Ulx5+iMQ/8nuBy5UJ8xRKZCSzioSj2uWzkhltZfaoFd8K2l5UB3rbBO
C3NEny9TVIIiaFCt7s+tBaWqoxtHcV/KukiJd/I5g3UjmD2NygawY9iD2dZwHLc1SyiNBudUATah
TyeHxBKHKgYirt7bN6sVMk/W/3LLkEb9N1kCigLVOkX68k7abrPrGyXqXpfkfq14OOdyCi+acLEn
1RWLys0L8UlJ0408N3INJ16EMdfXKFu0Jjisweco1O04maTRxkbLjQEuqAfQRW1gxGmeOkcZsW//
ciWvmHjjtBd45XTjLE/UubSjaQeRsR2m6xATKFDoB1HC33Qsm9FHiHmTPBObqx8C9DnKq3pIbJKm
PW+28S4/TUcNGp8zoCOK73fU5QGqUBkjvpR9GumPcuSszg8lYiUp/SxVtAA06xaifyJUzgWlh3Zf
LVAbPpRXTxVuQ1XjTVHcSUBIr4YhbXBuPQ8qtuao2rBbgAzBDw2E+GnnSR7tw8O8niZRNSEktK2r
4ETRvnNWMBOBF11OQCwbeoPTweR0aXOZw6wfPoEXBjX92pZyQd25r55YHnEuVW4FRdwO2+Wtzyls
0y3BvgoNm4NCLc5iNEjp63/NR32MotQFPrn0J8/vaO+650W5xcPAvIDWazyGnC5h9sJ8RHRUvTcL
SX0Vo+cHwNVwsCtEW+LqtzmiwhtO89TPkLiTGaQpjqNe9lYUS1+cKkE7QMA/w4qnnIcsnuOVDvCq
VCZUOuZqg0bdj6Hyu+9M2gBweTLEIYox0caL0mE/7aq298qMsNveEAz11ta3z1KbgpNTzv6bXPcp
0W4FN33X/Qt+MVy2eTj20L0Ps0653ZjOk2NiRGOwtwuRKbymH8IuVq/WABLYQGYKuwWbEzPzWmdU
aEseG4F4X65gEK7an9ExfctvLNkI4v2Bm5ITJ5lYZRuB67yHkwhIvGInGQBUVfNVjEOH2uoEx3dK
6pM+SGAimSw7gRFQTXuFudRsZWuM7dU18q257vxwA+rWMalHm+7izktuIgSr9+7fewrgmT9Ao7NW
d8uEAusmCVygoATo0D5IC/dPORwMJQk3do3trbaQWOwObhA3x0dxIJtR+z0FSWQTQBrFhNWddrmk
+OPjG/AT0xmfoaBeeJTXr733hpGMjy1OUka4cdurgedbTb+j2Db01vIZnb9yyfRHVLU/tla7ZR75
jctBv4poMq96oBzyST4EWzBrfxPZlhKtq+DnYhfXmTYA4I6u2lMO+U20k5EtfeRzQtvbZnFJcD/G
TCkIzY4H4crX0QgDxM+9gff4o77Glq/1i7SVouMD0Rebs37T6M5ZKsZO1yCyOocoj7q21HPYuvAh
923irE11LSArCpu6Uw33/aPjFHVy7mi8I0oeGq6WqiLM8AGurXYn8/8HgfbGNSF0LdMCXI+34S3d
XfKS40MEbOFeT+Hgnau7y0o+vBMhsc8R3CL5Ooz48tdUf8b7Hm3YzJjnXyFXIRN9Mg95bPCA6+N1
h4LNjkGd65uhPVBiqWG6VgZDzTjSIxHwjls7kTsDY3+oWIz5MhxnTRfExUOI1Qa+gMalK+4Dhmkd
eOB6mWDHL72zQC0AxiCUEZLe5XTOs8NvQRTpZIeXEWolBglV2zd0j4/aIJEX/qGqyworO7wwVDZi
lmjEhjwhiW1YIrmMoRFbUU2WZBaf86rEhYY+5e3WB52KF71nqLZ6/wjEPNilqwTTf8w0krJfapp+
bWFdHQA/g/PiLQxR7BxOmc32ayGarVOBP3bYZDRtK915Uj2xUoAOwIoe7iogH6ji8/bKkR9pOyn0
yWgSRomxo7bhSokKlb9CoqWFFYXiPdvXJQU82ehC6h4Y/QtjodTvXKyMQzh2T+mmfIteBUW/BCPK
wx+B3Gd6TyS7BWdVDDPt+2oMt/fLaF7WJaN6vfYj2r1uzjDIsmvNuR/CwaEHWb+KbTAwc8wyFGuk
bcDCWPrbImVTBxUNGkwvSeeOmPMKZG3fZinhff0k9uw3TqaDhgVQ/c1/4z968g6RhXrgFseWNlIQ
vWXZH7VA0j5LY8CA6k2HGa9SvT8J2lBHVaDJAaQyeS5eMDzUAZ/OS3e6HUCQQHjPh34jSZQDN5Ya
emgXKtpTNqdfZPZyUX841DxrYZEJ8rUlanHiR6xJI1xfaasZYcKvSAYwoApfU3GKmxzpUS1rGNZU
jENiCEMiDvPxMsdM9Ucq9EImIvy93XAHdFh7pdu/dtMfR1BrQWBA4M5f7pM3I2C9Hgz/SjDl4aV+
MN/muASrYWdqwKlbO/d14J+LuXKyxKp3Hfna5Rwc/fJY3sJjga8sRenjPTXJszHL58peBwYNQN9t
BhTf4w2Wbdf3KGrgJhEj/GZLqdpn78m1v39CBHtAHF5yEuBD+h+62STXD9N1cUdYINCHLJ9W2D0T
TGnQw+zuMKULfdOsVlTdHQqqDvQjVpZICbnjFrYzNgtEMk7UXFuW9gwz5OFRPTr+2yu3yyYhG19Z
CxTgYPyuTiMj5I51aw61PvZp6G6IxaOYv+XQzP0LPe7C9QZAgm8vYRb1jczGWHhuOFU2IioSBw/e
ifH4SSNZQK/80ZPqhuq/g0gtWECVRXt+PL6VyII1nVXR07jTStH6B/+7ey5owMl1yM50DwQFl1R+
K5fgDscd6m7xRRUEDrX/9r31QoeKwjV+4XB0wWTaoeC3tuSc43GrAJ0+RkXEi3SiHprjlF4P5mbO
M1qjLdfqN93BBuMAOqNHDU/WN4ettRBEFMtNkEJ9j3HCT6AnWOq4csTDdgQ0SjvsqYugVkpxbcCc
BHgsAp0zCoGjFEQnzyreM1kic6EZN70NfjzNWkG9WBwNHNyVWynGCijt26oLZQLzhRT67f6khbB7
6IHy4adYkzbhwxaXmBhc4BArNVQ+Z/OlHJW8POz9nSVFIum+aRUvi7D+OLsFU5SZ8uXGMmL2c8ZD
eBZxgaGj0oiW4DOCy3DS8LqbgIGCPnl4zh3wu8wKS2yTzQnJ9H9AT9ZgxSOituBtzpKKFz/KCQ5O
6g2PMANVut9vusqbqbmNZJWxtKDL7oVpwWt3MHGblyd/BwNOAsC1FA5Qcc2ZQMHXVex6gkYqqLwP
NpcqWNR3YNSGUFybAlpgAeg1eF2ip6IaRSj1fECI8J9xaC4/vxBgIkuxhgoesCrZo5SEhMTj4neG
TmishwIeleQmsK3u4s3En4JXImrI91tV8vZAp3+eqrGYofEpjW8HhBqHfEfl1b5f/OgATmotjX89
jaSMwtcxKzsO4xWreTfdp/hVNQ5ayClm79cMR9fcXIRMUTioXGqu+tfbUNF3JsOEp+gJFST/nGvp
dra2/y9Gq5X6SJdjGZe6ND5e49T+sJ4ayQHnG4H8/k9Xc5l7Xk5GszF/d5F/lZUQOAJxN/UBlYoL
j+Gu/BZiRpSPofIwUMw7ZfesNhnVlkDDOFySFcQpYfKN3xYvEPROhyrfl2vrl3m+QIa0MO/GFLzi
/kXFSmDY6FtkCeNl+iq7K1YUgtmR7v0+UDrZICfYOiIVeyEih8TBoKNBUTHL2k2EVu/41kXQ0Dg/
jRSp/QrhKg1BA/3EQlxCabnc7rJjD9RkEe2Pus8LGEK4wefIG3DO1Y3a9ovo1NiRXggBR9y6lL/S
GJ8CQn0ig6z6jLWioiYTfT5cjqZ7mEXW3UhRUuqfyjRxs8fqFWXh5dxlrIbNA1lou5yCxWavQ1sb
SNLMGTyxp3+CIc5JKv3sxI9fe1O/+lCZFHmIsuFoBsLK1IdtPKq07YHmI1v7r5uj+34Pmmk6S2Z+
WCC4GyE8w3LPiZejAcEXwMRXwbkKF5Hxz5jEGiNYQe5dfjSB97QEay9cHUgQFaB+XXZAxhs3Lq3h
lTls+2vS5jWkCX+AAEhcuRYdMwEUUMQ9iTnQLppG3oMV27pblAneiOp1d27YxVH8m3lL8OzooGC7
4CE25kq2lICOOpEq1+g0u7KQAvjmfZqxR9P1OfiYKaE4/ky7PzWSzYLYPeiUQIn0NGgqS80A6tju
HDsCdlqpY8QA4pvziAuOcxRGLHeav7jSaoDEJ+VjjdYUrPSp7SeaB5E0StwGcWXsEKX/BO36gW3G
UjtDpiYAts+8NI6lctxCyR/3ffMFhGZ68NTGDuKXLn5VtelQGaLg7nKRuqO+hTqzFT46ZfyN8vCd
axkwvBnjqnimkrTmzt+MpuW9VVp0Bu93INmVETI31Kl4fCwKegqMMlq9lMcOLmU9rGWhrQ5OjWsO
YsxmqeulNpoM1GNDSOY4uvbootftquKtK6ZtR+BvF2loUcJdoySeBohVqB0bu/YeTQWHPBKy1kdn
azhOiuv0uobC4NQjTFACUutJCDBP/z9p292ce6/fA3SclrikVajB9xBwzUjndnhVr6ILJYHkkqVi
uGMXcP+WKVnavxs+3hnX0UelhjHj4gwD1LW016T+V/3LkiMh3+6lueAGNNbkCo+3Jdu8+ndoud1u
Dk5iQP6SjEfgGLuVzTYZB1tbQqkzi7I25+8mBOulBQXpPMZTviku2Tf/woUJLY0JncYvC4HxQrR2
IIBI2s0FuP3wOU/fzbj2Nz8WOY6ThZIg6qQ9R3SEdSMpD+xFCdmb/Cfje0NDFZ/Qsbrs0ACIK3n3
wJQhDPfJIKWI/6ufoWKMj7IQqGUcEFvQVGxYcbhWHCv9gDI/w0rqdYsa3ipkCNG+lJ3NrIRtBCP/
Eavfh/ZXm2oKf+5FAijLmyPxdM5H9gTC5dWsqBJPqrpKPtQeNlm+NVyUuB6Ic/7hcnxxvmxpewtu
F7d4K59vmny9pn6GV0qdB/gSAjR1c1ld7uZwGRjODcmIQxVbKc1P0efbqrGZU1KUaJmCuo1qx5nN
Fivi1FH4VVW9FSgpDuZvetNwwNWFUU2Pi17bL2pYNSbacU7h5CwsZCs6/V5Xgv5scq8mi6vZZ6lw
90V5IVtVtUScVRFpLSsxjaIEQi40Fl1JrDhTcms9QJXNmZAg8CihfL1qtjbjIA210pgi9xxT+Msz
LeZ/AbpgfS/CrHRE1rpbV3L9uDX13ZGT7ohnbUEu5FtetElxEfCxtXns6jZl1dQ93vFMFitQgsDD
zAd7R8aE0iqRSUJA97hqIEm55jIVNQYzM+6hkjYuSVFcpajxj3qoec1Q20Zc9h2qD+nHZ+rb3g0Y
aKoUJV9TQb4PVUXW4m/wQqT09sPnf+JVV9dyfPPCBPNGtymhyIf0frAHzsLsbWasUlfUyCBpLJN5
CGjSbfTbm/PBdLx5A5SlEbb/hXSLE1yYO/QHWAjK7NzFiabOEb2huoDCQo00VAdHUlm6MaKAFvCd
/qB1Bm5lATbLxwVnXBDr8GFVJA3xMFZX56+BsgdfAmdAmW572PEuNu2k5DcDbZzQJLMcj8sQ9KFl
bT5+0JHPD3JknMz3dlI0W+C/PM0WcQB5/RuOe+Re2w9I07AxSocyZELFmyXipgsPRIAs7sv3DVuX
iNP3KQz6y85wE3ajAg2dum+t7nQqjSQ4ktl8XXd5ElLkjN7b8xoI3HQc5bW49rx3Y7vZOZGc+Hyf
qa1WzrKGopH9B3jhQIHYH7wenC2Nz8q1biFYPu2UOhqc6E1dWANeTjy0XayPeyAyvSZgyTEY6ld1
Jj4j3cuGJ4PL9jVY0oElKgOAvxCNbZKYwXG2y3adkqiv4/PLOGC73FE3bwo9wYxjSSlVvpkX/J0V
RVPXcTqFBhzHjQjSFdcmSteZAKL5VmglAext0P2ffU8tPvwyzS+KxZxexNOsvNGcWeNu6pNPFCih
hRZ7LEg2yg4wKLKqpF7Z4YVIIGU7rL6mjLeXSZ6yw5FGOkP7ia7fRYONKh/smZuhuyC5peWWyCqn
gUkNVOaQFbyruU26wgZxoFIDXW+FrLsYcQ1fIV8gzy8h+L2KAIRdepQ/5ZLQfAy+DYzQjNx3E0U+
wHSryHPbba8s3jXGZKoFTRkUBo1sx6PCbCWbpYKleFxBeF5mF1WqQz5OVt0fV8NKGU7QVh4qjsqi
Iebvoq6vGiXhYQFn27ZiS6AooELutS8QMgUDSBbKAsG5/x9rGpHagDF1WlSDvVKTd7oQW2DQkEH4
Xn2Q3cxgMPAoPma63H08GO6BH83Uo4yniOO6271BX0ywmnH1DG+ERf/imX/c+SiBf+iPFRgAgSuM
XS5nA/dhUoiinlbrDzZWe+FBUkGwckCrCa92gzZZSYlXBCW3sQpeP2DBd0FuSKF7sDux8hLbaZpe
VFm4CupYwaZg8MLivGTzXOxKbhbmDmlYFRbHK/wdgkbX08zGoJaX4oj2wcO+VZyDwEi0HTEqAavL
w73EyzRuuXUvrzJCqOPhat+H7+V9dxzh5bwl2ecmV28V/d8gNfSJWIFCRWCP8lPUInHVWI9qKWRH
RqyESLw1Zb76gPcciEmV9XrZ90litW+PAdsK7TGLWSgSIbFE34XwS6uBR9ns/cJD0k8uQ8JTD9Je
ssr8hlOExR9xhKNuW/7me2XOHI560Cjx5dewY+TWSw/c9Lq8w0y1Rp3sldmBXF7mpw4ujYrv8Mav
/bymigg3tUZKaoiVzhIxGDe812Knklo0dAXPc+I7FlOOwf1C8VVpxA2yZc1pRng3iVIlRhyM2wzN
udcf7GPfDLEMoZMOMTregLz6SmQD0zyLXXK0CK9bBfHzEfb3s/O2C6rLShZp65eHVQnuP28mEYhB
M5mjHUzDNqxyY0tSCqY6iLTlVNQeqTctw4WBdOqubKSxg7oO8dyy2UzA0jlmW3ZLacINZq2wNkpJ
ZkBQ1D8EmxExY1xxm42Hbu4v/OF1oTSe2XOwexXfs01h1QFtYy08aDFI0CQopd8fPN1eatWNWsUU
Ptu6WkzgSviQmL9aIWZSX/YA3EX1i3W9F8AlZW6mMBCTYBUoFSuRpplBOgM/RXVPsLOF9LBtgePu
reDdjRBk4QqVupKTlzxkq9LTUtn6aNu/lImtvIFfndofGow8wk5oJEOxlSe//oE1UymDJ/LOXBn4
GnLppub6dqFwX7/1PVd2jmJcTl9A8sokjtTGMkyv7Z6xaJpepfbWbUl5L71F5pPmyJlKO11Kg2Hw
MrDR3B7wGS2VnocjqjPYPNRYPtlgnweqmW1PrCFH6TzxoXGURQfAQMkUpNt1sOBNLGW1kBdWyzrU
PmrK8ssLb6DvwqRLxF/WvRm07mKz7t/uBWDD7dT0NHCnKmF/0q14k9kE4Z/Iisb1+PikGIGI9JI6
46LwUCd0blBxK8lQ4QhuAWfTXBhHMf92XIdgJj+mJZSL+yXieDyrpNAMFtgLpsqsZ0smca1BZbvy
uamoCt3vrQxK5NN1B2qz4GJ34rS+bDTSxe5JAXitMOdHMHu+3YqSSZIj2pcX69pisfGFODnBcakR
dZzghB2NhSb04L59jtQ+hntIhB1t6s98t37G7gzHq5jjE1Jiyxkxgemvaoue/RE57FmvMOYzCc2b
jOMZ4OdGXArKbbegn2VJP0ZfFrae2r9AMXLKSfdBRrMS/sxEv5eCwm7KeXoU+KC+4nV8T5Z6PB6T
OXo7GQueSPNV0D8t00OH2xLju96FiDXff0HXyZCtWpu8riCWIixH3NGQoM42n1wHjHO7dh0gH7yh
+zlJnYiSujHkOVeSZ2an+GeXVaputqy3nn441fkf3r3fN2pOJF223CzLv6IlPWtMAZvib3HXn75H
VQOs9dZtqzgr8QM2cmVerSfbZhNvkyfQU1f1d6lC12KnDz7CtH+8tKIw6A08Ww9XZ9R5N6zA3WpA
sdJ270aeQ4mKohU15CKSu//Ay3QLE7Cfn5Y+soRWAny6zbjur77H0eIiZ1rCYP2/AyfsjDuGTpmJ
qtqGJw6g8Olt+9ARLAkAnTFBW1mG8jgXzjhHLyeTAXJO4KjnGeG8WiyP8S9cqHK9fL8mTniHy75I
kU5ZcKdRwpcBV/hXz7tzUcNWnClTOyzvCxfIrg9aERbT7GuGohFMqvj3pPA8slLcC1QYm/WOiEqW
hDjZGTbNiUi+yVqQ0mITeYbD6hvS+D69wOpugPJy18eK0UPwdnHVJOrM1e4Kq6xvkRxeAZz6zY3f
ncNIwmHAD5i+GVjmA7Vfb+nEoTe8krAkWgXX243osYF0uzOxrCHubSV1rqBfrjIZXCh6qkJ+v0Bg
VXYpkZm7THDmTPFeKGEDeXNyq/Ssl4NWrY3RJosEzlzCVXb/O1qo/4AIbIqiWAgb4m9JPS1lUwzw
TMx4pAQCebtT+itLQMSA6fzgDjT8C9y97fw3RVonGN5Jh+fbXHprkMMtLeLt9Dn6b8UY9BfHp5Rd
YCgAhMYIZ6H8TOp7gcDL47DbYsH/ap6VpFy/xCNCkPBS6XUofFnGBta1AnZVNPfqYw8LK2TfMp/P
EJUpleotuxlPTUk9+8tRfkj1mpKsOKkR+7EG0RfttW53UbGUioioMUJsam3DjBZh4auHnxj7W23r
dXlVqhKB/7nuicBGsZOeR/NCrQTUi6ep0B1s4c4Y/YzCeLPOc+Rn1d1Zr+3QxEC7JVX1Z/ukCdEr
NLGEzOqGAEB2w51Bi6s2ZDubfwaR9C85F97FKvB/Vc1XJM5JAXw+d/yoXCIyeUJn6Y4+PVHdNvaC
9xAa5DdSgU6lhicaaq9XswPbog/CamTreqbhRWaRBJ/W0PD71S+vA15aTdQ70yh30LXgNN1EndfU
rqUVj6NpTtixWKIf8W1bt8AEk01KSLdhzpgZA2d3ypNn1+V6Q8Shpfey33pBqCQBNrERF9kGyJF4
96H29io4Z+6YbnnUJekC7+7xAHtBjFuOaLOnBrKKy0lXN2oETot3mMxDvRN5hKIRxSLWm2GkuLKJ
mqM4IjFtl50A2qsBde9tF9i7bkU75z5mmONtvnA71yrsw+/tUTbyf8xisKNcWj7BC6RdJ8uBb3IU
4H8i5XE997RluZ1MiDmoz9b9+XzP24do/UMVmCPtTkfsLn+gW2W3balAq0cefvvXvDmlt+ljlv5I
ATBqpflZqF9/3VtTNHZhHQNei1TBkZbR/og4k++ks5TEGl3TEaXeQmyKqWIhoNxdu+8nEtQ8UEdO
BA7ddHYyo47WdkEarWTkGVYD2g2BAtsx0SLDv7YBx6qlf5OvSLk5zYqsds7baZYXnQhGU9VWlT6V
X65iVvKPTXsjhQPqerQhMoigF0meBueYyRI+1f8OhiDQ7Gu6XY8/15P0glzAspvGhqQM2WGercam
11cAyPm4WoaKgZHLiZ7kIDAzBlKD52ZvE2W/SgZakjz90cHjk+zkR1acJ3/nosMGN/dG7ENp5L2/
A0dQona8FB8nLzguABaDw+EFh6HuYIxsb00+U0Kqc9PE7Okn01UlHMRlT4VaE422rLMFQ4CS14p4
jHC5DP90TCLaCzcswY0q5wzyjFkP44tUZfdmKKNGWz4iFyswIfA/6k6dm5c0beHUVfIJGMbb/u/e
yKCsSZacPbUNa1+QQdyBg5GAbMQLIjrpgs6LJBmTQMPNx9rk9sntxwpWZrC+J2ATgzNZkONiil/s
eG+L+Y71LEv9PxnLMrHTQBMj8nAwJ9AlW5ihvSCWIse0z88Ed6O9Pk9+Y+bJ/S5FWIWHo1cEZ8bP
wTVZolJkpZulIl2M2dOswIP381brwaZd5dr5CclozLpqFj1ilAD7N+trsK/p55oKaMeGN+J1lQqS
1XnIfvbY1OnUCkPdb648sLjRWZQDJdCaoSbyLgDGK8rPsAsJiEtZA+xavl4XmimDRnUSuO4DC5Dl
xjQeWWg8C/6XO3U051inL2/3zzRZfKlGkSeNsaaxlQO/qbuaYR9FRsHnjlTCKyRIv3OiAjrdFVqF
hReINRlqlUL6FivpB2v0D9w/zc01OX5V0Gsn9gOkb3gCxY0Lj27LJZRPG8pZ0Ro5lkA5Y+q/DbRm
KoRdfsIQ537MhMJWjPOnVHdMVvC6K+5phHVc6E+cR5Dm8+1/coNc/fmgv5fHgRh9JrySll564d3M
za7iBzXm4SBx3SWjxtwKS0PTBYYEz25Bl2KsIXz9FrQqxGClyAE1o9aNB+4EhXibviykDz7Ozjr5
CDkKeJ6k8pEdin4hQoNm2Pf39r+182gwW/pb9QUcUsKNZ5TEvxPsg7EjqhFYjf9HHcydA94KuZmp
ziFDTCoTRlP1XLeu0OIWD4TrRbjSljLC04DnsloO2xmyBqazX4wT7mQCtAQtghwBe16MymVe5E9h
KCxz2cYoxtAAtV8vSqMPaqocvdU8LZd/cPi/KgS8DjRIGZS4dvCOgo9RIjVVfVQiVzuqZOXC9Eux
Ks9CsiX6psDN+kcqlC1KkWgbgGOFkwZxhL7RmeU+d9H83N5iCRXK4lDcRn+w34/KWenClejiCf5u
LsR9AGZioTSVJenYhbpda3Dx4Zz4m07/YfyqDQ0FRMRjiKBiIoHnrWjtqoGSZBIY4T7q4cmoDGlV
q/BGLKgkN1g5uLpHubHWA2Uap+zjo8un21Efbwc3sRbBcHgGnE8oM85tNV/bwsWgQZOteuSYR70u
De4F/OdqVF6m5z4NtzOYkjbiZHHgXIjTKyKOPhGSUncRzrHrEX8Eh6miYJHHPOI/Ta4MErpPME4g
ERjS02BJUp5oUPGeKgxPdskXpJ14w4iwtBQD2RVNBOVKhkZXuf/Jj0Emy0AhOlTiiPGRyjDor6JC
2DvCyvVEwjJnUP2pOpSQqlXamacDuPAZfX7OMp67x0aSDRvI0xSdnCvDnP/JCs6ebem0wrwReCx0
nKMWDC2QQV5ibAR5sEUpAaNGHqcEfRAfRYlBYva86+WHK7EUEx4uHuMKBKdS4Mjbl8PXNKZhRqfk
Su9hra4WuM2uRWNqXpMHybviUMb+Z1Ec5TNFcohG0CUJSAlHPbdVr2fuCjTiLPK+Tb24m9R1hVme
ux7eyKDjNVw5Ta9w32APNNIC3t4m0b6IMPDIv9zRsZ9eOhz/t9oXgWjJLHcEzjVZYbG5cdUPZac3
tKv1TqbV/TUEf4aWRyNS41H/J78idDLeqABcgej367F+x/bliscIiPti29tpIVwBYuFet+3hBNOk
o0I+3VD0A52M7xjj9nmPPTuGv7zCczCWIkg3TCxGzpmLFeyG3tzb9m7qBMidXECakhjo2e33dJ0E
rHcWLiukxuXhKEIVZ676uWPxuOCFhEKupN0kfcahlwDb2JTY/XiMfAEazVfJ6CcDbnfYFSfs+y8c
kxFS68Vp8E4dG0pF9NLIi+LwSP3zLtcNYvgOx/Q0CSUV+XqGeMQET7zQIHK7LQIH7yI/5RuP7tkf
u255WnBE+npBA/oNFycSFiMullALYKJCz+ZxLyukGMRDuG8j4zzAdfNWkLUAzw1OJ+wQlYn78KCQ
n8SSoiAuSL0CAVt3IpdTk1ai8i4T9NHrobiVdB41qEJ96UIlGyiEqlKnMBnK/S4HO7hwgIRl+FPh
u6DDmx1iOdg9mxLjSsOF4kQtLd76MfXA4xuZJxtgmFkH5Ly//EUZdfa4RmNKjUPRh2KyP0KQ97v2
lOmPpDpGahDkeqPOzaggA1jHB1TigVZamwwZX0otP9PdLEnB14wDPgdxkyjgjE/9BaBrhuTPOXeM
Pswwh8a5qwqwqDRu4AwB+Jtqn2NJsICYn0kGMqMw/1+ochxf5UIPxK+EyN4nBkygxkFcy1IQj2q/
cf347zGbkg4J8u9Wje+b5SxLgB9fxVnkhnYlaHGyrwkEcgVvgCoONkAPiupXGTKaoK+mGJcRrxjr
02zDA1xfNX8Ggb2FEkQ2XsJAHD2vmY+YqiYtT6J+p10hOsyA6Rk9i//n6kn08Vc8c6BHydQDWRtS
zYOo6K9uDgq9AMqsLCDGZjF+i/bghwEQfz1727Bmuq88ZmXlCa+k5jR7lE8vPZrNFVzkWxWM/ygE
bOZfJFMTYFRTX3nNmTIkOoJknG5bcTu2m12fxm4PcV1mrs5X4zaeqI2FzHlHRIi0Xqvl8DS3JYPO
cHMkwqU5U/sxKLOD7YN5bl+7/PM+6yrU4pR4n42zdRApb4Tm+NKRESLJzstl8N8XD+zOSfv830kz
jurTOutNI3JHL0V4Xv4otMbh8amVTaio+FMrIFlbHi6m4Nc+bFQOaMqPWiSClkzCq3bXEERf6Bq5
8jvwPkBRy9t5KavCOauLHEOmNXDJhC9ABJN+ZTUtaWJV3emlYz64PsHv1eHykkRdmmWjE52iYTiS
U1f11qAJliEpLnHl+E0ujbJQ5nEro3PCsUNmlfI4wNx8enj96EAAUYm26qbvLGRzRMypSjIlVPTV
v19NYQt299ER9cKId1KMyzG+e1PXklPOmTjm4tlhLSOcN2qorfZvXBtfA+Js0IoVC8OUB2JORHHN
cABJO/WwAgqXFgvwUC+W+x90i74n4HGfPPge3yYY34ReIPUDgMwbhmVu8zPu/4srl5Ax22r3MXOx
HBWRjoyGDw8sqMBbOyH7VtAg3N0OPm6XUlWHBiAGime6jcRvitPHuDZRPD9ETMqUfjE+ClXYAADj
oMsuGIpeaUxqdGtvLYVKd69mYdaNobbwpIqo2MnwbkWHTgOvJ0jfYpjKaPVrYGnG8r0tLz3lvc49
bSNlocRW+VStc9EjaoHdHOz6BAdLSu75FUVuG8HGw30uH5Wm7PFdAsKNy3TbB2zSPduVy2681FHu
z1d2aClvlhBwZiJFZBCNeJjaNI1IsRTf0CEfXwrlX+j1Io5cO46hUfdOGk+f4icvlReuSPIjurua
3yEfYIjhkCuH7YBTiGZliZ/+nbsfY6lLHOyt7a2BWS4p6OoaKHIq+DVfJ5GTMuA4tuWaQqxEaFMz
MFpJRAaZEK71J/t2v9gwXGNlXBpObRqoyPV1CBgJuAF3Yo5LRDCeUT+4IALOnVwSvID0MaplWAiX
jOxIgnLw9/fko1eFPZrxCPllEzccWsRtvtaf+qalPqwuBOTDyDU3tbEO+Riq4Y8Ywi+/nibXOyFh
XRlzoJT2EwBuF/9I61AxBiCxQLi+K6KzLpQLGBk3RI6bfUMD1Sq1J18NKHuBi7wB42Kl59KCLSR+
VB9psdKrLM2RraHgUsqzGcP7lT92f4zGE28JVvKVFFfNyUfvoB1SFy7+TGnqoG8fXex7j9y+9AMm
syQH290eCNTTF3xrjvu3CYQBreOq9dCJ11zeW+D3vfuGk6Df6bKRS+vsIiH6c+3fV8DXA61c/zGm
xe7TtyLBFe469/vE+H/Zw+GXl2UHSK159yWxx1Ur8ZruqkZjBAF5RABYLygpy62yqNYd4ysp8NwF
iUVWqEjKgBPsrOlFSBTqKhxviAABiPlfCdP0bXA1i9uakckCR8asCB3LSUUf1w3/703jeJCA79YX
VRE14xTx30HQ+RNQsuZe+29CfPEZKHPw2iQgvbDL/C3Z4cgJuT3x3csIPhM+R6bveBM0oU70x5/e
CTvtG4BJdcNH2zmjqM3Uk7IncduNCwuFXky+l1cWGtNpulePVXilF+3mCszY/ToHabtALdNPKuKe
1EeovqGROxO+ESo5gHtRK7ezYVfiG0xRtuvb9Ldgk7OJ3s6Mw641MatBnGKXinJlKmL9GH6nJSey
Id3zDng02RVI2/HZXUnS10re+gx54o0OsuJz50V+VCsPsdrW7vTCQy+2QuZpKO7n7CAoqp6sPHlU
YsXpez28rUJlCrUAEEWS+YAB9/tbDJFpGdGclLxeb/P3uRdSTI7O85Ic0lGjLGPdGxnTJaLq2ro4
Eo9JZHSJ2LYKJIYoxeWxKAu5T2vPFwqwyEccuF7apd273uTCjDUSaZ+kwXIe/ZOjVr6f5CAagwMG
5JmAbaVFJrYEfkAobjPObgA2ADC1Z+3jZdaWtm8PW9ijQ1Ad+pS05UIO1icsoEzZGRoWKPDJ6wKL
re0JijUO8AoIofaozLV/7zUl1gt9KTr9/ErQfr+I8d/NoOJUYMoc6gSwVpfH/U6bPqhOi3R4Y/jf
7EuUZO1cucBo8wV8IM04PNvDsZY00sZYgI6QTjmx0/Q17uURtDMTPgpWmNICLnKHonCnSh2sji0t
f4dPOWDuAzxLIw/+2DxWYTtR92q044SXZmhl5OaiR2NNGUq084+eZS3W4hT3IcxaJXV9AlWUHijy
pMS6Vj6svdYkTUBYLtiMCEDKwlZjIbkLeNXFqjMvVec9gsL0tSEAUgAirpCMC+t5akpMPNAalBqa
FsrKy6uf40Nu1c8VSgfIwaBeUVnKmuLtD1wvoYU4o6NT4kvBzTtmGOJMRqsiSS1g+ftN/12RqONa
xMDZBHuZhpOABph+NEhPz5eWu0l+iFCuE7NwUSkc0KW0vQFDORO9ig/nCjTg3vKvIgXmx7f2y0dh
0iervMeO3VH4NWnpcgzehbJ4E7aOTRpn+Z/J7Y++BepAPVlU9V6l+fl+HPW0eugKgt3LbIavlUqg
q8uP+sR8lXoGaA3cnfdZH67xbjVdCkPhjKTF5dQCltnZ3fALIu/2kiWfD9sP/Z1eIaIWHjz0ghFr
wLPGrwswItUyd6hdUfX6RP7QO4dXlu/Ji60zdz/uCpLMXAAyonSKbYWL94jy+9OkwKe567gjW+GO
em9sTFzt2wROlCKLN/uoLDiQHNkPYlGDJN4I7vg1lblZSffQ1j/kdJ2eO+qKJeLmA1VR53oP+40E
bLlSLFEG83atxF7Fd9/UWwgtEz4mDtWq2yzTpnpFZ/ZFdMWg7hZsDx4OD6qP/i7OJDUjU/ApLR2S
Glu6dYeknLDZYW8XsPUfjRv9PjRvyDl4jfdefyC1CLPz3To7jx34ADFmf/aN519A7ZeTqN+QaFLq
kHPYs/anN56h85NgNjKNrq4tOlOhmj9pxvEg6KZk9mkyVhbJtgmK90ZQv7K7AqYYD65LSWxIap2N
Y5RSf4nqWKvOFjqR4cAv9kaxmNET0wkIDcW6oSHY9QZGCbx037jEYd1+z/26kyGYRtPraXLTRl+h
kFNOk3cLRH2cecJ7CIpbtYI/0HnMG4u7x5lcvaqPKy0kjXm/KmnQoTv07jvUcNFNnsWEjilUl/7A
7l+VQ5YTjxDj87NqnQUHdVewozG9cRl9tjFSQqWeweibiU9mf3dPMrMB9UoKxq1T5WfPJ+2UTGb9
OeOyLT/wzYE25LKVoYDJwzCPpS7ARGJHe6EEUXIA8mySHFbO4N8+6yV0KjjSlhczB9jUP4Zt1Dfs
Vx8I1FujoIFElHHFZCr4Xlc7IqoSRCXHDzCnt26l5PGus4KohwrtaOHlIf5X4SbvhHcJIUHgJAz6
7+oYo+1/HLg4tOIyjzTD5Arv991deIxucfFIIE94NC6cZxPCV+qqPlasnrpwoVM7Am1cIUos7ET+
6GsUBbmyPrmwjgtttJPtdZcuourtaegmFuHvW2zp9iNdA0jIkUTg7ZKaW9blzzKsFbZZXc7AhzuA
L5YM1LIK7mh/uq/K+VeobgPCtmdQtOI/WQoi/XmiIu86ofe5+UUeKiv5e4jNIHXtSs2J3TyOXSEw
+0YtLe7Pp6Ek3BWsfkX7QymAB6LP50QRHPqNfJM2AJxZZPfGFmS0F7rItMWK9iZvJmlgWeZ8/vok
js03ZqjpAxDnbUS3evWnZLBb6dGLyusAusK/Jplp12ndmObUAYbCJMSA80qX/qQ3aI5e+MDhELSY
RgTLeDHOGcTYgk98lJIV6V+cBRXg5V09Nyind5pMoUMSxrr7jhydIYPwwDCNRyp5j/HL3ATDmqci
lyEZg69qttOnuSG8fu5qnGbnjU0UpzSrfhsgQt9jJTgpULS7Lx2TBd2Z/uQemabB8Tn5UVwaLRan
x8UsetxP4efeA1QHL8pBVT2lscN1RigTRY88Sy3dwdp+8gqtRaMcsKm1YrqOqY07RV7hBwUuR9XM
CnApd3ULhSet06h8vkPWX2AuVaPr7f+/+gs64SfoS3hUeqn4o/kasc4rKI8e+bBbR9GjNBfHA32W
vLKs+66qAQit5rLns8kfPLWtd2NuZONh/D2MEXziQERi1zcRbxvnXTHhNZXjfcZK9XNS3FfTa1iN
yqUVsKpb8fSZcwU8cZ7lAXorJjioWr/VSgvzpOXXlG5FU4oQk5DeBJENyfsRgHEnm7yLLhPNMQVz
NYkD63So8uqvujBVI6rWBflNNAe11/u9YsBDGmYG6rIM9hXQnEOVuOCXHWqLaNTsbf2Vb4ixbdsq
ZmzCKOO6Z4BN1pFrtTlX9hsZfag/AWBj0JODPzj62vqtg2s0bB8OBkhbfZhAPmCkoOsGoKhzz1ue
P1oz4oDdK+Pv/J9W5EtUSsNZ1FD+KIJPQ07PvYveeowKZzNTQ9hFRzHjx9fYQrQtMHThP1+M1GyT
R/njTwzwCdvJj2Z/NvgIFQ/FqIWKekciYAprhbXCVIoGZ55kwpJNWqs1YeZFofSjiSPTyME9D7xO
FWy6EAv8Xno6aDIT39LrB2KV/D3CexH/tl/dbgX5z11E8Lm74y25I+5B9xMkEJbIGRYo/98azdtX
JNyI8MJLqUhowWyGY9ktd8FxAZAXuoHiughptH88HX/E2hCGFHDTsRzhH09GktkjSpQMdnEEW41P
OC7EEoMxCWYlvbDeSFx0AZF0Y8VWbJbDFNjlO4w6UQVycye0GSrNCTaiWHwEeo9/4nhqc+j1EFoA
yFY1KYhubYMWeZsln6q/uPq9f0JraMG6R75YQwVTMYd4LIVNDNwDf4OWgm7Y0fVraYkPLwaG/r7o
jhlMgUwklNMAbqtuwH3ixnWFlCbFBN20eIHz2hch4J28n3VsbhlVWqxUYVA0GTHF+ZrUmuedZHjA
/GWd/k7BfmpuREcrV5ztXCSU5TDxjezHSVZJyQi7TLhCrnnejfRVkXDwOxPHKxGoRsJq4mCjHuKY
1FcLmV4BDC/DrcXhJTGyki8U9BDQTYig+CWr0BmRF5CR9PtISTCzveE/AuTraSwdU8GNVAyRWz48
go7rd0kjitx0xRLKQCc18KDenTrSHp830YtV3lD0KV32gUkISk3WC4nB7S4SsI4M59nyNde7FSUx
cpi/qfcBCnWGGZ9GndV4WJyR6Z8GzQR0tSUkYWzpX98fGX7YtjTryHkay452oopwKr19LcQ5NXzq
u8J3AEfu/u96mXRM0G5pRRw4y3M9LNNn63YOwb551pMm/D3iHK/6t9lubEkanunP5ERgsWgrFt6B
8KkB+jH80AWhvmaq4Xsv91A5TXSmsAETsM8D8q/AisiGpRcEt67jcw+htRdYDWIGF2rq0Dbnt0mo
7ovC3ecE0SP5A6ZwBf8QkWmf0aS0Hn7zQl2fSDB1/yHHaw3zLjISScke4/Y5kcYDqdqM4asCI+6H
jLcnOMsH7oOjo9AznPpacQgUnL/iM75vK9Jtm6DlZ2uoz80qS0WUxv1t46yDZ+3lUiNTAtb55qWB
URDbgFBnFsyqI79QbLTbwfcRWNdCtMKvxfKCGc0JaX4bZCdg+USCE8YdV0YuWxIzV/uqQrjWBJO9
/rDeoDhAZ4SZv17CrSIbDPpP0Zq3Ao7dW9N1g+7grJEzBHTgiDFeWJnaNYygIFpfE6vh/Ue5pRQZ
eUx74mW6s8Sgf1SV8dhmRtp8TKZ6CbBXbAKRTbbJcwHICExHFamQ3xBY5coUZIrC8fKswy/va7fz
KNJYU2Qe3SFWInHnxVg90r9eUbvz++cZI54bRua+2iFQtPWkhIw9Iyh8WfiO91UmGB32pN7i3Iee
rbPfgat8brPDVS9kSbI4WhAmF4u50bDI81eaTc9fuxYpELVZO3aPmxBoK9AJ7+A/+94fTINTYJpl
+HC4QaK2DGmUSZ8c4hT8QXzFdSVq66JBUrEe9KcSxRb5zXQSTDCkQk2rJojmKqv2r/anQLH+yzcw
9ZZby7Z1OmDLtwzqGoHfrRgLvVBpRfMvei4yfnzpt3Zu/I2Bpkgoj5BZTDCIKL6vP8sDrFkjgIER
3aCmg7RZapElEFMQ2lbo4bsED0Ch5pvKaGmwn0tAv5rXrJXvEdAMHy4NBH1Az6kcmtlE4w1yCa4v
Q32mek6HbrsWMLLoTxbdpgfldbEQIWK9AA06ETCOAZhylFYlf+OfaawOJMghsMjHsFtasgT/ukSq
Agn4XvZzn1kWNQt29IrXlH001PHeiKQ1H1yTtBAygnRi+hHTlDTl5x4O4TT8TaJVmCai0MTSE4Xx
detrVzUSIRLVc3neL6LyD0ZtCcarw37GC8whDKLfM9Y5bSC40m/ccgr/BQOUvGSsNKo/rugcRAWg
W+QKAhIqhk+kFiJBGmm6dtGn/zaZYD7EfoNiDFAgu6FonheEHSaHsRtEmN0ux7awwcTyyLghsM1L
1Av+wS/pwH2JNY5aUs2qnbfntOcnDXUKAD4thxet6PunWpX6r/NDL3RCnHiMmaZ0OBziWQoUyZ97
Z9wtTFr1VW235KPgCN5946UJt46NuVUnO/LKsthdgABpMmubhhwy49TeQPpZ6u6GkV6AtuXtO6tj
uLdnDefz9nHwu14g+VnmnwcTU1zLkQSSIjRrTs6UI2jk3dUNrkaXDllXD012eTht4JQVpjEq5NF2
qI3ywkS9O9nkxczwOEXS8+h1UrmzC7DvQgmzJL3sKPr5t9fQQ3xQHo1AaaIJpDqjCbcI+fcbkUOI
JqThfDeAhjEQc0H3yy7XWnmf+Sn8nKuInBwCTCPCynYRxT8hnUDK/aVXSx6FOJYkmkLONSQrjwoq
3uvuROgeYjKLy8e7Ky7S57BAsNLLV6Cr/0wtoy8fZhh6GhHjM14WZnbxmi6SBMeYk2/3zJ+GR6tU
dcEKwkzlnnvRmFnJYQfl7tL6K+2NiD8f+uXWKw+xTIaFJ/mBHW8Nuoak1yAoPxHoJLSh4057C8D/
jqeyt6nceJvcwNroPemrS5jvP1JFnkdQaKLQSLla9421XBjDC/ikZ24kbia9TohSmkJ1Do4A7RoA
jjaVfklpTuQEk0wrirKDVuJ38b02q+HZZtYVQ2Q8/6g2keWQOaeTlPsdhxJmerxcH/cZRNT9API/
4c77+tTc/keBBESTh68LbNAuI1b8I2OAKo1+wlkjNSyiKpGSfC99AW8z9eIF1GXbiH5d7Om3a/m1
7LVaQvMN+smBmR6eZ04uGl5klswCCyFl33aixdeWXklLVObQXf12Hri/YqrkMFmtsCP5hFusix9Z
aEZ/Kw9MGzKEevDpSgkGnzlYTc1mf3bvxeLmcfI6F47S9mWo3kM8zb8dZJ+lyo3TqiQrGS+4Ot0L
hi6S3wA+9plTyeoR2G/EBqOmg/HcyxSkYYWxggw8U35pHfJU15e9jax7rHBr80a0BWiQyctmjupX
N8Qh0iI46hc815hbqxWYeKoxAAKfDkBv+7KXvGG84z5iO+zAMgRB/TM6o8CMSYqRMGu55745GCdY
AFWaNezOL+1Z4uNaV6UrNzxru/n3HLhrHz/mVuY3W3UEXKOmPIS4qBc9xmbcfbnO17NjlRYQ/QXL
sn4sVTleeCNBIs5QVmc5zTYiUve58UfgcXFJAKnGoLpcqIC8+rJvb1vR3VMwsHDwPdlHNU95sUJW
MiEuSI+GYpVvZ18/fJma+F2ML2SMKcIKB9sBDleWAEYDQzo550SPuPdLm2mDKEEb7ibfCXZMgrZa
Hn+k5wsz2KZU7wNGxevnGdhzqV/1Ql1Z28tsC+FIrUt7rF4ZhqRDPD7EysntS/e9GN2vbXolKGhV
MRAfh9udWcqE/8iN+Ev3XjIb4N8ewmXOVgRZA/VFfScKnxflGDe+gz2IDQyWENZWtlslqeIjpqzM
LjGuyrYckGI1WYby+tBdvxNuAhkC1cMuwuGGPE/IGoKU1W/jJI9gCh+g6EAQ01py//CjNzZWkVS3
04Fnf9BF1JtNAmHXi6jxSpfJl9glO+TY0/iSTWTkU//ZZoUro/PVMQwFZOLz5Z2Ws78yVshaCtk8
Jpcm6boqK+fWrkvnfxpLBZpmpG6Q5lssII5GXGGeFUd7J2h+x1qZa9XJv1N3Il53y4oMj1cSv0P8
yq1NduLqB4K1A3afbvZhpYN8/k1hvwM1u91JNPhxItub++O0Vnym1tq6wJkcZ0CKdvq9s7rH0p+N
Rq3JFiLoAqoOGlFarYc0SbLJZGoyBeq276GKFnCqoksVZ4jyKF2uKD9eCs4ZmG/bMFyfASUU0/xO
zgtSB17KzsqC77oNuzKemv8SO61ATphyJQ1NB8y6oKHBmpbRMs174x/mhZHxvnvOrEfitmaL1uwN
zZxKrcHhcc7tDN6HwExQmSjfgSe/3ckOP3NNg1QpavNhkNVlqMB02Tv5MmrtZD4pF8cttDnbZIR0
orO2I1lvwJQiQYLcf/lv8ttaV3FLmSEdxQhiU42hpTN4h61DZiygywfDfzWY7CNAn6k4okxyoVYt
W6sYJ69BqbjblkLIhBVInfzTTElPZen02UquANt/bkFszbLbJc27+QNclQHsH8kLGYHXv9xjnmUM
A2AzooSQIvd9aU3E/FaAOqBD5+cfWJQjwIFcQ17QJropCIyBqh/BfXy1SwC7VbSd1gj7I9jruGk4
BaFk6LMrTnfaYDD44mIJrSXqwDYKbl6RwoPXhG/QQ8cZBCvhtqwLlB4l02JjbUN8jjNuSh2qiDRR
aeXyhDsh4V73/c+pRkBl2sad1MP74wFDd8KjSKBvfYQkxqfARbBo3x26vwVXllJraTHq9tNZHQ0n
Py4vw6JkHpK7l/9RU/wR7GbeOG58k9WNDuYU9h7+SHvFS06ah3m3qYWsmAUJls+OxPDIDfOxwOka
AvHbyr3LnrM35ubyr24AfRTs7MLXTXcnNt3cdDt0tI+0xspO7uWoIGuH98msfRcpywyv9GG7240i
ldcXJIRoIpzeZ4HQ8ovhl8qKUSdwtcSwhGCGMSzlgteTRPsls8eHlsrYDHxftH6fkZr2oFpn3NcQ
ridtJ8oEsiR/JZ9x82YPlxwJiQDRs/ti7J603lEdxJfI3qC+4ZnRHmEx3dp2dKF03rnOUNQojfHx
JqOz+Jm72TyZgWT5BQDZNh8MIJzKUXwhUUwHr0gntM96ZZ9NQ9PKI/aowKckxvOMpdqIvVMy0NdZ
E3/rZwF3WaCI981Vfso81ou+C5kYUQIPPhnmL8KHs1PePNT9YiGvivSiUx36/KCiPr1IPFqbkDj6
sUQML8lhYgSrXYDyISM+14GY0JscyP3H1ZBdav8cLGfFLjIKWlefNIV/UG8zWvoUjUFJmQ8m30jo
iLEupcQFuOxRON0Avrc1VKLqIQ33/Ts0r8q3l3+Qf+bl7XOJqciykyK2vhzuTLna34054QPWR8n4
ONgFUx1CuFo1lA3Ooqg013wr828xoyUZI+nGwca9uJi8+NTPJgTCTzEGUUhEEH13AilFNYv4utKt
1wUoSTJpNG6OlWyHAyfkonWHSSCHw1REs3O4u07v8FA0C22IPnh3s9hdKKKlmdUDtCKzc65foqfn
ugO06baQr5uhX48mFkxkWVpl/AVJAdl9sMu8UXwaDpS0zf7xdfa00EN4RL+DWaKd4zmx20nea4FH
XG1mQyWpewVtIKp7576l6EB4v/NsEKJdmouTU5A6fXs+iv2ed15dT8M/dLG0hSyoQdEP0GynugJx
rAaRE38fbeVdfpts/tlIUX/jzn+hKUuzqTSXNCf+NWB63WhV+HoHxIThEOIE0qMmnpBZ1K46GHgE
MXxn1NDFgX2ktAnwxdiIFMYmGT1XWy2GV2bxPHMV33FQhKql1MoXHoKjlUGTwEgCjdDby1I/xVyz
xproi1yrsOG4OOllvAozknRdZHYzcvA5p8xVJ1U7i69asbnsUWX+rp3OL8zuG9bZ0E3tcMuG34K+
JfTvE3keCTm/FY0EosxublqkyTzJYd7JNI7xWFNjbTlvvVrCtzdfBT58spnQQElKYKcFD0ElPu9u
HO8Rq9WfM2rfzU4ph368nUGpNaGiGAM0i+yvVO6Lx/fn5EjRv3LqWhVlyQVLNmKlevhj3PVljCrO
SSx1Uxj6Fm2w93jX57M9JuL87oZEH1zA6allObvaGB2pwdZoh9CbW5VBl+PHNYaJfNnYg8bj+dsU
S8Fkl1Oq6JhnFlhD56MKKXJjaOkHPn+fne6tiOfaN9PG5/8JAlEpdjorIQVkRdtSSepVxXYesLro
bSh31LX54JInVKNJD/Q5oAsO3+slSGEnXSbr3392Ja7xf5MUaaRSiYUqPI935HFFkx4L4plIHaRF
mi57nkLhusRfsUr5WVJmcGeotcE1N9jeMSzkgcY2rCj3sFWOEYj65XmYK1Xr7ilVJN9O/x1c9kYt
DVdSXvGioZvGa7m/yMx2pvr1H73Pxp7cx+UDlnFJb5jiJklljS7k3q5VPZJjiI671OGrjqkQ8huZ
WCZDMlVRVw8DG6TjIQk8Squmu+hrydB83Ma29k4tUqSFBbh1W8JqW/6jNnnXuqGDzArBd+c8yDX3
getkjYa+QnlvIztjHeYUURhW7LYP0pvzh8yMXFKIScuXRoGj5Nf3qQttsFFHiMRzl2sNEzwyvHxT
fFH6HwO6tq/bcW0kwSuyT6wqF2qoSG29ayxsS68QFjk2dcOkC6S18qxbo9qtW88cnVlqbgxauCYH
byGQxQiAIsjKfBteXzEemUz1ctX0FCEFZy6pxm4sgtpHTFcj/Vfb5YxcXNja5CIIL6b2kgP9lb5w
pmbGBIde+NluubF/Ka9AUkuLr7zP71PcbZUJdGbXqeYIQDX/sBwBLI2/6n+NUdr/8PGiJL75Raqr
kDl6I8sAfd9b3M25FmDzPsbNAwHlKaApCy9Eb0kVrMXvtKvcuY6rCyXCbJoLFSbhRUMIPeCF7g4p
+fGHAfp+LWJ3FT8DDiCQ0YPdthyd2QxJNAJ9sg7Z8q/4R6DXemUmANeuGeOUXJWCh+Wj6irQpKW2
3Rn8iu6w/wEqn3I/V+b+8idzq3/nAi1G1FLFVxItOlcXTml+CFWQsNSHD0qf0Wa/PSunX+kIn6XX
5NhI6gN7xF1Y1w8cXbK/m+dD34XmCqeJuBxVDgIjFQG6AL45VkWAkH0MaPfPzIGw8rNu8oF4zaRA
9PBsOBnn/nNXaAxQckW0Bwk91o0/HkGpikSDwM2ZCMs0NZ7IgxpM/VEHkP0do1KwAXTVaTafNaPi
rsgm5J5XCeqA6l1T49C+wZexTmb52wvoTj+jhlCOhaDY1deV2iafmAA3cJrUlnt7DVNYm5+Sr8v8
54JcxO8A09yXm819FOM7AkkZJJHFC14zfl6XuTq+gAQrSeBIFLpLBOEalYdz9kxb4V0w8nTVqWc+
KE9JoZinc1nlHZxcee6OD/zuVpgCn880ruZ5Ru4hDk30Dsm2VbffiM18P1ElMcCbYgrD2AmMB365
2fuJlYxvsf2kIS1Lxt6CQN1Mm0Ya6f78fQhMRT/emtULY4pAptoy2udSp5vmAglnlaB1p6faMQwE
5I7Ydf6drIgNQ+aGTYGkEMWBD5AmC8D3gA/Rcax5LXxfNQmw0q1gAkL52J20NVMoNcvBrOINQbNo
rI1h5BakvcWu7YGUivYNxSLcO9ZmpS8fpK+5hfWngESSq9PFrJxyfpQLRICoP2pdE4XC47brPDhj
gUQgI/yvFqUWJAnlBJDu2biUKtzC/0yiiC8ErXEeOyjgAgw7/3IeSmBfoBUHLwwgwJj7UuOK7925
oUE10pXpxvAnYGC13KQt/ZxDGKofTYwd8i5S2wXYRqBxt/21EI8vnFbiZK8KgEjoyKFkwnob/x5h
RNFpmNYMGJ2iyvkisALYkbfCijJDSvxuhPts7mFaokH6ihmn3HtxKhSIjkvMoewdD3Qv4uW4rbXW
y02sRKlhWUb9FuoQpUOojLfB/SrfFlW9KTz9cfXEzsCYiqP0WJ3LuwM5UNQ4zSZqoN3qGeGnWcze
G9C1o/LRHrR5CocciX6QKwzhiyQftcfOToHol0SaqseAZjSbOXUzADJQlvu0ZtkMHiqazUpwQLK5
Rsv/9BzRqboZ300a3/rrF3uh6uyepY9mtpmQAH7lCS7JMpWh8fn3xhlUmFHqjCTtS+Cl0zoHQg0i
FhwQGr4xOGusGyKQK+4X4o/j7L3mqmeAnqLzw1wkv4RCREhjUpE+24Jd0NJ0t1I0VnUDVSwkZ7Dm
dOttf/5Ev6oh8QKJPbrsicLI05ZBtVsZqVEzrl4m3VA7MVYOaraGavZLxHuaW/7EsJOqy9QlAIHc
8SZDIKdZOzAG/MCM417BebcqlvvnQ1vgFMU3/Wqak0s2lUjGDUGLrp39KI80wE91lrKQHGoYoBYR
MR9+MFQL8iVORbv7arGrigV1OkaePDE7Wfas6b66IvWoeV9VaaS9VBl7IhDZsYzk46FPhkPMi6gS
Jfvpn3GqSSbaPUeI5GC3SLN6FU6BFt63ATwLTd71FVSQiy4vgHQOMX2qyi4K7CIFZKYMpPzJxZXM
Gu+Mizhffp71AQ2b5cW/Kv1Z6xmMAL3DqSio/hbuwykBLdkXk+KCo+hxRtOdxVImHTRBEs90W2/K
DfdtO/5Q8YioBzijXQcK12ieAPttLr0FT1vQJ98TfBfVYOq843ydBRbsCS2OM/lzIc6OWRfz6MZF
C7yJQNAQTO+/6MHLm3VSFb9LvIgtGprdoxEHdP7vQgzp19rNq6EuSrRtpLh0sopngVZm5723PvBh
VvVikskMzLwJrPzr2LW03hQohrCvTpcK7RwuKG9339waRClkGKFnFI4jfrgbSRzPtWk49CwOMxji
DzixED2rK8HIK54a5cixITEGkclkzifmZ6U6P6Y0fMD/Zst8g4AMdInnCOwkKqKYmySj1GRL0yNQ
2lSpt9hd47nqt+vgb2WZmxpCJQeIbmgGgm2kz2gPa6rABlHaPM7EquMzZbdU/og4TXQxGESJddXy
tUgoD/Zyksy7OJWOurPjfSYmUENXhuvZrlU87pLOl2C8EONfaVM8I+MwJEv+AiWfojsb/oI0X2Rs
874x98xUyM73oTURD2EeasFiZFHfd5IxNMMYfWKqEZJoKri5giZZ4jAEVnLPmtumFIG4knAEVSJi
uoPucIiBMD+uSEwgLJG3SSBMvfK5F2JrTB4lw8EWaaFqO7LtYHPekU1foesVAtTcU+79mwk2331F
gbmmzehtzTrkelrgvy0FMc3BUflxzucqkeWTqYL96Rw3sXanvxLMIOdXrHXnDHE9XSUyJUpmOhD8
81NbNnlloc2jBkgN0X885h2XThKXXoqSycKUSYcS5g8xuoGfoe1ceKhR7NV3p+BnSYIv05iutP90
nCyOErw23uGXApgC2cskGECJ8D3vbc/DfmR1LwzylMz2AqcIXedvShJc0P6imMSZoFyphE8frxys
ZKsk1eEVUW60loHzAlLB/IMWpbkE+PWrVXWalXLAwCQD00ZUDSuWfFZuaqvYto/k8v5IkKm11ZnV
isD1m+cWLYm3spkhp+lmDpkzeU3SO/MD8ZGrRcVfirSexoi7ey00N3uSf9lsyeB8wjudwDVYP5Dn
Fs3sRVsSpL4FCfECZp/Jhiu5/gN/tyhpVuK9U2HSTaaHSTdhtPoS9JEq5rXIStJMZsQa4nfBrN8T
4qX85OSfwUXjTkx42o53rJffSrUxM/oXQBWEe+Azzlah5INzX1zOUECD+M2+FEw9/Z6RsdP9hU65
qz6xGNFvhbJXPaefjfmfG7XcqSlWEVETi5a4ZTy+Df3rdk41hD1memOzPZgADdPG0/CvyLl4isQH
HMyET/0gFdlsFnEzJAkedia1xJ/2jzuy7RtIGRf/zwitkgQ1q7ShNBZB2aZ981XRBMYepAIR0zyp
CZrf64EpbUjdfN+7dP3DDEpa5dlX9C3/KjsxxOFxkivxRy0+pDvNm39li7y3b4V5yvq7QgF0WCil
yOy3NRlTuIxSMRsWaO1jNVM0kjZ34wwjV594z+wuEDGTJAQTF4KGK/PaY9Xaxarnb7aGa72bBnIe
2ZAXrOCm02qYec1lhZLOdvS94l6WWEPGvjgnPzHeKw/caQyncrJCLF8Rikeom8Sr5zrw8AB9sPD4
vDEjdh0wOhFnQt/9Gtv7n4lW3PFI4iWLYBUQMphc/eFad8fPqYp54dlkJC2sXOxXpvyzJV/3Kr/y
lahKu1mc45i7KEG7L0NGodIflfxugrJ6vkeuvDVBXJueKKYkRUz1sHTTuWsfrseBdVzLCPmQC66z
/I/bfKXX1kVXKOF2hy0ILNWHKuFbofVH8/2n8Qpe6DVwnJujyZtI7woGmLdeGtgTDBCmGg0TvOoQ
PV3FwB9VDw0M6+JtUk3UzvhJyEtxQZc9NthsK1Xt9cIF4PFwnfs0tOYMSzBHJYqqs9oNTaPAmRw6
/9ZnZxebLcd1NC+UK2crei3EocBlzF2e6AnbGuEzIzvk620JxYtEHTcjJ8A5HfQsn67MoIIygxZd
jblnTLO+jb7FULF0zke5G6yBU1GWPYWhUhaU4jCjtlhczspl5Cq21FWbDWrwfkWHU6aRQiHcTU9h
C1m9d6UTb29n3gB0F3xQSCMnNqHyCKGCQvQtlKVX8KUf/Qenp2YGP1DNN/S1A33q7o6bWIJ9yZqB
uZmzn6xKcw7JxTLRQ3KzRV0UUZASTPFZNOVclBRa7a4U6Noc+65LQYsjQnkt3DfrMJbUXMrWd9RA
WyqyqzUIg882guli31w+YYO9eWepD3HEvArBsBoCc74+3V5tr7lZIjXADlCwSYoLOLPMj8PYiTss
UDQrwOLjZl72XwcLuGSp2VNlnGJNdUKlvdnDdZ9ozhVZoJ/Lc7kwyctkdeO3Pcj7IGHDSj+cUXY7
pjSJI0G+lz7o9xBu7vnZQW5a+FfifGcy8H5jwyjnQxYUmnWikfpmA89yvSxo3Esf2yrgTyBSQSWA
DZUargl5hqKWHJDkGesWekkkBtMWbYkexY/i8LN7FgEofHYiKeMz1IHAqLeYse7BzjwVCF7Bxw/3
wQe4v0SYBhgdUfNxvn8e9aVCgbg/lh7H2oggVI+lvMdIiwl6ntuShFl+9yHk6AMkITC+ZAUDZ5Ab
IPEQPN54OYbQ/f+2b7O4u08DGuUOIsDfeXz+JJuD89eEi7NO1joSJIyG+jo/9V2v9j/aePVJxes9
CJk0ap44tCdKoSRefzHjBW1YRyOf4qLIY+hT/H3g9pAl82rNhPSkJN6ecpFzd4dxddPWs/z4Ge0i
J6btfRl69kjQpQzkEbWpV+Ed7CqACTKu9oZbyLfXnfjxvf+VPpRTi7+JqoJ0DF9en/+DWK4+xWVE
Busion6Ck9RyzS325rrHiSINQHE5VWzsU3xzi00/GQVOmWh+3rF+FUB3xvPuv5dqXsBfT8on4T22
kO9raObN8fyEXcub3e8Cv1KoJPpsUht9x+pJ7BEHQS5wQzpTcTEMGDYEqV4plrlEswSkRHL/XQvY
r9UR9q9EVYujZM81+mYyFkLODETJvIqHDHbalydp9Gk18F4ElzmmDGU66nZE9d/2hZDP4VbcJh0j
ukWneL+C05dYTv2jvQd8RIywqlQ7h6QGRqypfq4qK9Mrf+pltvzYvALoqiizdkLt6BCC87ewVMqu
SqXAARwoJIdlpgwZo3CUdj+ip2W86G5pMuJJcJ0litJhwLCN/jENJ8GOVofr/t5LUky6kGBrdAgC
+5UOPmceFUS0e7+TNB9z0Olxlae649Xt1LhGNMaFOeQ5UbOjTxGT2x/BGiQCr8VP1HhQRBeprpvb
oMNEdbXk5CkHm8CqMJ1W5aVfCTJFn8c3X7TdjltofUGR3f6uuzTlJfWJyebFhOQDriYN5PlkVqXD
ohLqRqmExcGpOPcAwFNoPMo/fslpBj0q9SczIGCpxzYhF4Zv89pxwJkOICRDcHJINF6ySxhDb818
L5qV+gHhXdLSnPKOH1qisJeaxeF0+gdVTYqR4QIoxlMSHkYHBYJRFJTvzIK/1D+bd2tXaAlYhCNh
L9ADw1aw8AxE+SnuxfiR+Rh8gwj7gqZfHOHofb5XkcgRAKFKOzqm1BGCmlx4A6TQzesyaQIWNO9X
WyBh4CtUcPEvzvHVVb6/fajuaehajRxfINJQ+/HMVrGoFtPUcsRLt5wD6sx2ayNtcUk2DAevb8+C
GRMZy6ITXwJUiGhNhoHdYDi8a6LJgZemZm8ETN1Ax+fJUZ0YHd7wA7Kr+mWlryfw77IBpS1L41KM
9DXSuPxj92vJTDxp+0Pj71pUJRfGv3GPvNk4KKiQ1iyXnNjzCWGYtryt2xmFxVvwyCrU55RLCVn6
2ODdJ2hrhjNi1mfv01bOtMwPkoLJJuXgfzoLEFmeojNbniiSIa7GUnAgE0Lx4cO6aRdjHqY7y1o5
DYYdD2ulZ4P4lR0z2wa1ChQ3HDFGyvXZqrTAx9FAaP2Do1YbJ4N67nZk75ZL/MzsMcB2VBYqkP/Q
bJj/kRzDc6o7YCUETW5/Il2LD4EgMfolkb6M8hFQVvnjwyBEI5etizgU9C8VZwTgb2ifNzdS2fk+
R2tpD7u10Viejx2+TxOgzpRixDgBxccV7iPfNewJdSJ7cmxYhPMDs9A8cMT6Rp3BuzsVAPGcQqEo
rUwra3d45p9j9siYdLbfuXQEQm56r6FcxUm9/9mTcW/rLffk2Js77f2ncTlUwfeKINf7tyIdfTCl
/U9Z4DE9hs6hzn8SmAZMPkisvN/+By3S+xnZ3i/80fINcYFaymC26fnjkDZRiZqPUca9cumbGtBW
hU6aW4vCvvbFis6Xbawivj7Rg+OjD+JvIPru7DQ4QzJSu4VVJrkMxQX4Be0yX00Vbw1Ab45nxiQE
ltQ7FyGimJKbaCvL7AaKPj+/2zrEF1VbeHsmGt4MDiBlImOwH62N5QbRlXXAtFvAVpIvAwnq2doT
U5x4F6VD9gatUWiSzedNoTPAtgE9DyreSS7IfJrUZD3XozWALvWQT2nX8KByxd8AiYP/Zk5tPaSd
40fTSZRNipzUemlmPOLlThb2v1R6uXq9QqnZ4KbtQGSGEuZewuURT7dKDxjIfLVTrZ71umEEHABt
4PIIVVQTGKKI9tm+EIq4ctNIM+5aY8kqd2iCUKNiW3V8jkgkzzAWY3bXUDTaAa/MLHCf/Ps0miZT
ndvj7PBSpytEoVRk3W6XfB6BHud6y2g5WGaLtcttx8g29CKlpfYNDGXNIC916mPxGW0DFRhgQtyI
Z0LLcuEMZZA8eGQvSrNbhycuggFURZcuGTc0PYIRaZDjVyUw0DYM+vFBYDxf+fuNrh6lQRMgJBhP
f3ecejnwm61cO1dFQrUawbarJRJguH1pOabT8GDtXw6x3AR8t4ozohxLJHfVrWqadqpf4aYP+IK7
blrVZExkfgK3GF6nrPEDiMQ9sJfbGzp4g5pV/i5m4voPQZ5cQaxmTJOrs7ehQqiNghLcWLKkFGXw
xCnTn/Ez9ISj6e3zOizPVajVolzWc1xEmYpCrvH2n7jDdxRMvuZfymmzRVYBedzl1+a8qoRwtmsc
SbitM9Zaar7+Gd5NdDd+Mh7d3u6U2vwWLXW3O436W2qeWTuh+DT7eB4l2213c1OaQ/DodfVoftVV
5euxtCYuQAF3cERAxcEK3Edd+a1jVdVaOgofctysttGE7hWlgCH69X2jFp0FtsobohK7e1Nf+CJi
VedvfUAc7Clt/+F/QuhUboZdg5jYZ01AMl3tl9pUDKoYEh7Wbfpjhmh5n8PzucleZHjcKKBDBfAR
9dlcINCeobjy2e6rYRvBSge0vR+4ri0cXS691WhPizLNYGkJOCR4nkcX89sipgleSFLFSZXpPecm
aYxZi3EPXhZiHJpkRgN9gezHlfAk6Bx/GWIXckVHLY/TX4vqj3vUCrVFHcjHUyITCz3P6hGtXRRA
lDPUGS4qdg7Ad5liLXUOribqC5tOSO61eW48bF3xrbz2X6iJ6rMPZPSDd/QSEC19vOLAEYnx6UGO
F0A6VRcwWsTkaG6PNac7fttdvunn+uSx1eckVzzwNP6wFUhxLLsIASotCLjzDQpw1DbVNcjfHNsq
XdWShQSKe4v9kYU7Cn4My3ifJbnfryg6YrK4r8/fyDKFzt6dhac5VVblIuDfTXJSy5UYY9WMtmFK
G87rIykPWDgL3KLRzHQ5yyphH7a4cZUYTnenMufMood44OvZbIJ7YBsoIV2J8akR268g6GYyO77e
OmKr58JvWWDigsZH4l8jogoWzzRrpx9GBZFM40wiznHLYqWl9m0+Rw0sF4ajfGiIO2810MU8Cf+g
1NquwyUFtlFPJvFovKqcfUDdcHfHPpE8ANbP+4FWGjF7rmbnTciD7g3ckfuC9EpE6mxJUh2hH165
3IhrdmBUdxC2tNZue91rcq4m4vFhu//Z7d1MI1MbtD5I/zaa+f7V24jiFHRyMkxUXEhNWkJlpRCR
y1YeBekHA37xvwCFQPQSBiV5PQeROQ76zJF9DVV8nh9T8qOL9XJHeKceiqB8t12/LYY1Lh4X71cZ
YblK21X5bbAHrnxc3XjljcWgDHna/lBhkbvkUN/ziZsMGWcWj4AZNG09eZzukzRlSwInTIUHAISA
9CHVNp6+COcz4zlQEnC4YH45i0drzZbmAASNLacHMHoA7Y4pEckHNQK0kFvYMTOSm4CymF/U29qJ
IC9D8LEjsaEPVmuOTqpSiEHZCvxRWokiXncaHez5jReGvvFsYHJvLnEE3rpgzvcQLQmNn2JwiK8i
W5cm30k19I96/KmDp7Y2t0DTxe4NJEOwxhrxWcNYD8TKs+hEhHvHWdIpyssFw81zElQjOLXdtACR
+cxM4vV/njpupgnOV/hcmlUbl9/Qy0/MzatwRtbD0D2Nr1fj4N50K83Sj+4me3bKMcU4f/Q6/Rfx
H57+lXh8kk1YEggGaNJ4lNUq+Xdf7Fc02mvT5UwGSb7/I4FfCnIVavYSmvJrBgQgDDJbJMVnCT6u
fb0OkQY0w3NIeziLhE398Cj3URFGDYuEVVt8puqxbxJfl9sjjWucq1Mru6jyv170ViQL/QRC9r7a
pC6GMaMZu6uN2PpxAPM8N6EuQhXivQU1XhNUZ9k3ME5872VBOB0GtQzoJJ26GxD2krEkf3IpR/4I
TKeQFPhVn6YBeuIV286TOzvmhFxuUaVdxq/TzBJB8xX6OmmoWQZvxnT9F+Fy5WR1wVmAYGBz0VS1
u9/pik5tc1q5JQbZDJoOf7xWzGtme2YPWaZEXNwXsULQsLST4j/ZrSJKGjQeGiLfTJVoaVcNhQux
prq7LEj3q7sEzDjueZoj8W5DrB9m1hwKd1uGN8M1uhebXhZ1pO38aSj33JwFs1NtcSxCR/UE/YzW
JbRMmPq2S4iSJ1j0GoAl6lUlo+WLyiqxjszCEXze+PcU78F8EYyXs+ijLSxCnFoebjwWCHjFC20h
8SCcORE99o06hPLyYmX+JaqDhEyB/sM9WYq4zBbhgy/6gP86hcoExCsG7qV/48e2mUN7gaOaEJ4l
WGBAMaGoVkEGdNJrnwZUjUmehtI0UsbP1Kcu4aIrpwkkRfHEySRPa3+OMDQ1sHnRRmvPdQcCWnW/
04i0eRUpJW4GwsR0Z5baAqcdvm698B8Mqyc0L9zoqB/SIYvAixYYtE9bGKBAtIPT0ntyhRXLHHrd
LZDaJi1sh2Wx5iepAIGHdWSIfeE8B1YddxsQHk2fXFGZLCy2B3Jdtt73HxD+hvq3UJsgb3bUjCP4
rQPBPN++Z8S7k1EpPaBlIfjQPxioPdMYlOGbFOyaHOQRySISj5vA7xKah9pJkxRXkf+5LNUT8eQM
G+LdNi3daVcDOWnhlImRawAzZOXazrjYgey+XCerUTaZvHstzEh3z+cdIaS1wfEw5jrvmyHT4yW5
gwWSFZwwz9UxvzKVCAWPAefzeMe0z+R9oFo+5nNZX9jhBN4g4fR2//FzJfQbSNFQDH4fEj4nGOQe
f8ZvTS0GnQAzFSdYVaZvJCUIzOV6hy2KA/dYdBWMQJYNLAMkSGAYmuxDuDuHXn+7XtK5f1Xf68zp
KsK5z+MkYqlCs19xKTfcNkMgxxR4Z86LTdtrgqaE69A9zZ9WjyTK3Jvomgi4T8u+sHPIwKZaa2e8
bpUIr0kDpOJK5PBODLTa6KJlZsqe+1T82/mCY/ivc5GXOsRLaA1gIzIs7pXMV8xrsWkUkTAuPVGm
9iZqhLt/VvAPj8O/ERupQxxp8+ZGHr+vGTpcPxokY1dMLkgyq/gfc4zVQ47OBM0desEDr/vdwNZb
us+2eVx+Fvzm93zZOuu8vvameQF32+nmPnvqA7haLFK7COhkDJDMbwh+vXt6tuZ9QwCFn1OTkpcE
wr27InEuYyMTHVnyd2lKyshQbWSaz7id42VR09jlXvza8FV6RNrT9krosat44vx0/Jl2G2/6QcP6
mw0ua1MC2/Ak56GxhL1BwaYy4kt8W0SJUEUygLHBoRxjJ8gOoewMQW5AdScZVzVX/mFmJUfBSQil
7uY4Kkgq6CeVyc/fTsY/7O0Ur7S9N2hVJn9R2+0S6tjBJq8EOgOQQwoHhwUbVzwIoRgHDTwKgErV
P7yRFKvGKuspt3DjqE5XHzuYs9kQqt3nFrrikzMlTPJd7z4KWWhppg/IQj/gPVMRUmgROVAdn3FZ
GnRo9qGdNrq64A5p8elVPNf28NstZXRZGINNIhUnO2D/ZMOyijJSGAL6F5jBKUTLZke6jwkfXadV
Wu6OurRR8HNhj31tzLQcoNMI/sQfg/VGtqLNswgyRBj729S1M8nkGaJs4LeFli+NtKNWmiJ+Djy3
24yinYSkgNVLT6KIx1rYwg0NmN04+CbT2v3KgiRt9BEB0AGgT7ao0xWjCkbjWbYBuMIHNHs+eZri
ed/WCw8CoG/nlsP3Pr/+CG2QuucdwqRQ1lyEj+1QO7/fPMo/97KXp9fh6heBqNQBD0VN5wWlqRKr
0GwPcRtkjBa66JsnRwx6ao7oIjlShtCgVm6fWsB8m62cbEqCb98Fw3OZq2FzaqwJvwsHK92cWPuw
7MY1tK106a5SudB3Ar/Wkzx4Ecl/4DQpZO/c14VhIWwOTfhWJxO69X6sIG7eSuz8V6f20PRC9zP7
1psefJP+6130z6KT4xhT+daktIz42o8FARl5Iu7tTBQmFK0L3/uBnzxS8IioKcCiLVDMnkWFBogt
6EFn7fMFAhPrKxEgFgu3Ii6SDZBa6X9Jm0y0i/J0VnK3kVLv95aED9HZzSPjNUXT1h2rSWK9aQ5G
Dc02XIyWkcuW7B/Le2g/pKbhFokFbCTKHloGPmrb6k1qg0ndxH1G6zG/WtQGSmFKvuAUyWRV/9iC
j5GVTStA6zsXtJZZlKFCyaJRR3Hlkb8U1iwNivr97HdQEQ7vtKHpI6oE2DJ+FAAVP8KuKO2z1aUc
DOO+f0CwLOaKZz0IQ24NcLK1PFZiHvRBfKTMD7Tsr6EYERB8dE0hi7OrmbMvP2LJjsOQG2IK9aW9
SfZu+mKYu0Km4ge1l4BVKnFaCFpsNDSm4gLoj1r5UwSzoUZDLftx8QxFnay5fSyp6dYofUUi7OmM
DzLGG1yrqNi245dg1wKXRmhWO5hb/yksoTPbFc2yKdwVEZ63DoT1u/ifa3mxh/usDEiVCzOaF+Qx
FDk2VTjrKc55MbYmZnVSRybWv8NJiQtCnpAQdUCjB2bWQITr+7ULJI3V9GzjaGwSsm89P2WN7pga
Ai/NuImUfvKsFoZYQV8C+lrDzLxXZw+pfN+79A07HIEZmDoGia4WPfsDfdISxlegPX60NzG1v7Oh
UPQ+bHhBXe6zbuwyHwdVx9o2HADggiV3HZOmEL2wTkhbzs+9Zgp3835jo4Me1cMV0krur4MQoZGU
l5Tv9ZTUOUV5b3FZWlQAqNFOdnCPk37BXthglzGB7W2Je/cIF54HkFU7wZD/1fnfZ9O6gADMovAH
C/8TPZJznm5zQvYeBiXEiKcA4NN83zVBw9aCHEh5JRdZmy8L+1pZBNpmS5sDQaMR3eGFUCR6tlWb
dwH/AUOzWrUPZjob6IPmYcwY7oWQ1NJItsqOdBHRsm0/3pcrTfbOC54UhUfskwBsiJBza4QZVHY8
qvBcLqpFOSQIe1q66DoqWwwcf851COspmBnpoWtbXJyxYRy7blEggStLcue0U1zo2NuvGfal6dQU
9/pYq8bdjEUC8HRvv+Gni3F9FyElwzarlexVUMnnSVCiQu4AjaH1BK+wHwjBy5B47BPaPx4eNAn/
mBsBCBRoKMi73scWsjXyie/xoMsbQwtRsaHO/ZKQ/+ehcXHvMzCoKAJv/lK5nJFqvJu7oxsBN3wm
ff57JGaL8856uhVh+Cq0PKvmut4UCfJM7OE2bYi8FLKk+NmQlnDCM6QcSfap7M0V3HFk5Ki6pmLR
rfEE0JjLHBQrkoMUVZeLlYzNtXwzRocv2ox9oRusZ4k/rYtQNrtGG4r/003P28Wi6PULmVa3zBaZ
NV0APGruKAukcDIu9o9K4E8QeGAZMISur8jDe5R6sLMlFPC2SGiyjXSlqJ9CEFHwwL+TJCXcEjwc
/lqeEMPs2up3eDozHOJB5zmg3NjypzxJ0YL4k5tNgFtAZFCk14yFpkk6IO3jgDij9mcZUdj76uaf
kHvcWKWwF3zPol4FleqbJpwJeksdDzukUHGdYBKQTOVKN36sVwyBH2RdFatiavkUjX0rkkJ8tLEm
bAKp3avZKNCR1PWe0MNC7P6JHMU4OWPk7yYkpVHgneR7t7XRrcoFo5S7Gb8HZEHqIubSCyQQd2jC
8stgzk45FBseoD6qX44tPQo1/naKm+ei7hrOD2hkh9N+L5aGFA3jldkS3mXhpbog831Hkb4QCYxK
+MSIdod/YS9+FUhDf1sr/VOWiU4++Z+7XNaawfX1wNbod41TdgCPezkRZwBiVhiCWP5jI1Eu0sEr
YU3xdjdGTMWFJI4j0WHCGOSOOt2aez44zhgz/xWpCLoklzOkicpJqu2qH69uz2ugYmVU4GMAmCZp
vIFbHAcJ4QwYfx3he629RPhs1WFAtZgg4blwShMnUT1LEgxbfmk3PXftqI+g/AOgoHxrVFCFeHLe
Q1oCZP3F2C6dknpd0VnS52ryetFAUGikXly2cM/CrfBMsNw3Ad628Zo/QKnXaYEkWzTm5AZTMPr2
6M9pV6jOzzqxDTIH4p7FRlEDAtTLOTz/oXRqwaqEOobO8RH2Jboox49Iz/jG6c7r+t9Xuf42oKf1
fS6RuHZwqo04/zCSIQ7mbVxhRjRh1PcAW6Tca17aojrFhnRlygdYyO8KAlpmptCMPOFq/9GXiELS
ubrgsBWOIi7ymQYm7LZ2HMl6ieAYvMx4q/W67azAzbRfddJ1GA3997bgwJiJ7QW0Cpv4TFG86a2K
a2BOd8+TxB0B5zQPPxgibUPu4p1QL0EpSZHQHUr+CuS+b77AEGDiScY/WjywDKl4dXcvQdMbOXZw
TIcuTyYuvZyr21g8aCAsQepM5fKXn9sbcm2L7SRFRvw1kqc7QVHWFGX/Sxsar/iWL4C7nmn9hUf+
8b2fcdfg4z1lTDwT2cJPsgRLQQbpHBEr/mWA0xHG2M6DsHLQ1YVGFOEL6hqKkXr4OxKkc0uQEKU9
nhx3OCCI1yTDKxVye2TnXM6TRdbRkgjwciQw+XFH0Jjv2sPAqW2qqU2/B5Gi9WZJTzkK2v4jLZdO
pV2z554osvSf0pruUCZgeJOfIVLDZSCLewjYBc4duHK3DwyyOMZuqMuIdQUstL9vFUvB62MF1AB3
u/Dx5tsmiOjnNTtMrW+e5qY4U15IO/dQve6e0OI0vw8pzkD84t6sBOCLaQTBDkpjmhwGQuWAEZeK
kZsHL6hUvHGypnUb6l44V4rJpUxNLe0S/sC/K1cQgEVcOUFAcASaNBI6MmSOqFMG8kYscxoX3efy
g2uKmEVA0+PzLRl3riAMxy5HR3dh0pimmV5ft9yzMmvNpJYO1gWg9mvzBeOAu9ww6l77iJqBvitq
vAUPi0zrU/CORzYMfaFqhEV41rDS10p4k8LKxj7EEqp5l6mvJcfl2Vn457XS2S2YAdXAX3j+p4Cz
xfNyFvzbs1jvC7dmdn49z6XK3UBV5rZtof6vedKct3qdSMrfRR2Im9bdB8Zu9STpCccp84BAN8wq
Sn2z/6rhg9FqrCCM9MoNoL3+1QpZ98AAzFE6qf+/z4V70U1xUIJ3nqWzdHa5GMo0k47W9Jeztk6Z
dj4fcXjXYoDr5yA4Hn5NAJKwkzv7yNOFFDX+MpDC/SjDN6mVoy6IQvZMulGwSGqIYjNetsKY6FP/
+Elq7lsCcd9fyPywWZOQsB9cjPWi6/ONHR9UXND7z2dyi0rMJnRp1of+vlZGtt06qfIWoAWGUNoB
dsjlb8cdW8KR2SKz4m/t55tfNOWrnaV37N6KDt+ct3oISLIwvWwjEFnATVgIO7zvijhcFRa0NOio
j+H0w22aslEmd2DuEq/lgRypSdBmh+yRp5lTGQBOyx16PS0WlBSRYew9q3GRnSXMoARYbkczJft2
tR4ab7+8EzC4NsDZRDFGq0SK7uxpgZWJWpYuCYB6TQEcQCqpI/KpeuSwZpsIJ/sC3hxdgOtG38GZ
AtyryHbO7trEbK/VgJ3cq12y3JvOQhoVKje57JpV0h/pBVmfR4J7JpRG6GGtLkhkhcHw4Szc7l3b
uZM4Usdo1WFGcRyIdisIK7VYUMcKul7WTcMtyjyf4tUx3f5X/te0ABqr+Ewk/DFDDoqLju+NAwKQ
LBcZNgZut/ZJebo6zvJtAaPZAnww9Zaf1oSuCOASmN2KfXRE3jmmTZb4i8ErdGZAG+3Au3LC97rm
aLhLSmJ/NRi5qGQzl84UjYGvxCbueMS2sFjv4whQzLKUHDrfJKvZlNxdXwmoMGWs9n6O8GWtxMR4
ZcFxR1WbmOIf5QpE+IKZlY9jZ/p5/GB6/CnG/BGqe0nepWQsj4JYUOOL0OU+iPnDPvPXP5yiAs3n
qQDqBiCEb/dnqhOvmPWSoSwG1V2Fh8ZBlTWrwAjNzZf3oViZfHv8IJ49WHza/LrB6ColSnoNDqOh
CkQExNwkEuXkGcmnWs+dfd/yTgkl8ApXgepKmFrhwT0100TgPpCjiTClMM/evGrUH7KOwtO+W0Oo
LWnLg5lnp9lxoXnohcI/4tUSYpKikXJ9m6O66Jt3PnuKZSx3nFjO3SfBw8pZdSGiah7tplCc9jAs
eM5iQTfeyfiggk6+krf2vcgrqLqzuCZCIkrL4FBV7RvyWhmSgYYL+flsufQaGeO9bLSQDdSlAWdr
0Z3WrvD1LD0qMP/F69iHkE+XauhfRz5nI/IV59AoEDqY+q45HkP5yS3RvgOyx3Jvz4MYemFWcXyT
E0+PLFbQFImoD4UZrRnR31ZxCImZw80GV6Yes65Qrlb5NPXdBZ18o7xJRdqVOhOGHFXorJ6s/tKN
abzf0Mg0DtCsp8etihXJX/FfYS5OjldfqcXVOoUqybkDQuXpzEkvrkJ96hrzQgCzKUpqJCbg1xKb
qL80GC+Wd6/WKri7HJTkt0AfVocvNKFJJqtNuA1GoRAVvFyuihfFb0azAXJyls03a++aEi5Cg5V7
y/4pj0jVFjEmatS4gbDrkinj+HFgRzy/l0lMUS1BRKg8PQIGeZHiF20SegIh0dDafY3jVUDwAwkI
shvp+1zAOql/AkdxxNoSaNaUUZ9h2wEckJ4PG7b7b2jW3iPPzEpsFx3Eb2mxDMtHYEY11I0AG2wd
4m+PX4fNI7f3e1807O2EDrUcMYTiEKUgBtt8v6uOevlkmUb8CWYGJaysrsYlaW0mOa3ifZ5+17y6
r//bZsnznb6erelrboMApu3tirf2Na9NiGlwu8LUxI0rzlF/B2eUeOlSQlpZR77iQnb9/aK3LFlV
9/Nq9Gdl4hheatd2dc76udh+Xif8kg6YyEYebzNp/guEQR9UEUi3gUtm7HPe5GZpROETeIcJIKGK
+44Znby9PEZBKkEUP/r70OGe2TQZefVffKQWX3fa9I/4Ii5lvWgTgP/cwAgLh4vahnSaKFX2raJb
lQvb9kYTnH1TfAFAz1aQjT5qGu5zgK1hcU3jAty9DA8CrA0XURDRrwOfnWMvByj/BZfvMEnkek4h
Cv1Xk0D5SQoamRRa6SUKL2fO1nBzaqlzQC6EfzEY8lwvqG4sO2rPQ8WCnNsRRNwhu7mep6xBezWA
ajBGVdhFoQ7P9xm+Vz+MZsjZefN3ROOrhRIjUF9ic8EMqmoYDqTySLVRH8SfSQGOYnJzkRTz3Czh
ofBzQyLau60uhIegG4loeXogH6GPzT0Jbar8CiIcKXekxmDAVTolrjXU47F69adHPjAI2+xBHIW9
L2mVKNNCe8qRWA5tANY8F4cHqAGLdqHBATOI0nKKO0sS3FdVauwtq/n7crVVOJfCTDmnneVx81Bq
2PcHxvJNh8RmZi3UL2/KNzoU6MkXZYBBXrmXEJX95drs95slCUbMshA2IWE6YXftTVCtDtWc+Qk6
zkxArr+1XX+9PUD0rVMhwTseTO/p+jIlVzAAg8MRWKDRjTAJ1Gs7SU5amG/EcfT9cFw7jY8Sg9sL
7MABjZ4EZJW3g4WSOVst1LX1VkhLq8BMJNx6AltnKs3WHeEE2djrK15wOtCx2t/uXLSITN1eatSq
z2QFNodHUr5bmNjrqT6wXumsUuiPCh6xzfsAJApMT4p4NGNzRxFbmo4KBmbHtP1XOIBdsRQWkVlH
x3O8cCHKq3wBHLmbbB/AZ8wH6mAAV+IE03/AfC5hF4iVdp0E1tVKzMh1dD2XF+0GrK1CpLVXZsOm
IWjn2hhYbmILaOr8w8wn5GRsvVzCTJEQUyNqfx4nMA6/wPqLInQWyN8k37slAiEzPr8CH/FMlIdA
ACjgbdGQ8jo1ytnkMyu9c6DmxEhEBzSjDC/mF0jbRMwgZTanyNOnmjghWmcdcrdopTkdMhgOM5Og
Tmp+VJSLAdKg7leuXYXBumaf1pEtEwyCpW9oCrtkXLNLP8p2LqdH+3LwaIQ9xaWHym/V0ZyERoWV
JpAd35xPxNqiGV4XUyYynZ3a5wVTgFq6lufukY5hM2zP6AWFDL0C6mWFqphZAAgpyfUCf40eeUMP
+jdTJVB9W4dPNOdkQrP+y0I90VDr+Skl5Icul+UG/RK/BOSbU9Oaioyt9ZUOvHpOMT3WewEn8CBS
6EoTs/JtOU1/+DOTsBa6i3eToACnOFNHGD9qDFJJym4vrXYGwg51kU6OGpumn0C3AaU5/Gb9SY8P
NWOBxgSsXeWGAAkEk/8q1UU9z7SLV09hFX3TdeLHCPCuwApv5lRbrtMhW+zLZsgJns0ck+M/3Wae
cFphzwro6Z/PAv2YvphrNwr27QAlomXjb3ScsUuRmsFm/YzCTOe0O7TiI8l/NAUrOuZZ4sZyj1Go
upU2lWx2FZAEk+Y3u8uOCYEhe/mVrjVsmewANRD61cj67wrCPLJuyNRFSCQ1xiUGwqLc9JjYlxhd
hJo2t1StL2uDzyg29emzixVN6drKaiTbOTUPHGSVbRNbxN4nKnMHLbBSvcG6Oyym7ndb+JoE/so4
y6utlMaogWZb6LeMmwllSu+3IrnxKwPNnmgfaXYHNU1unueQPQfXF7ok6vGuG8yllCUbIvwy7vP0
Bx2smWjlSHQ6aYi1EWd5bK50tgFve+5MOrpFSoDzbXFLQnegezGDzCmhbScc+xaM0RcRipi3smNL
+AylH81FvR/l+VGor1+wgCIrLfXyl2LeGaYQc/IcbU2RbfO+tcfVkKitiVAYxnMrzjCKgRbnAhfI
4+vnA9I8JK8AgkDfJlO0tn0fuQvZRQM4WawJMwQi7T3csDJZJVES8PrPeR5QuoBHFa99bJkdI7Fr
KHJ+PGb9R2u0ZLJtucNj6G6bTyMcaI8llGBdWTLq/8fnseUM4aSSoVZa2iysDk0+MkuBAxgSkdU4
XXUG9l+pdA8oX+x/VEZDjdcQcHMiBp55BqNkmd0GLXsZ64A2VmxgRxf4XYNFfaVagvbbUzygVCyA
FkyZ4o8Hxvz79Qfrzn6gDbzKG/hs2ViUj8TT2TXr6s0Bs5opJLeSZIzj1UGS4q1VuEb27A20KS7y
gDphsX8Uj9Fim8iUar8gUl0F/arjzVh5PQ+TgOFtBsSkNd/dI2A9MbTxy8NpkVGExzh65m5ZGgL4
6wXl1z1VsUzyseXIreCbcaOI3/mUEk4spVn0TUGP/KVYaObhQpnkTd8msoFfhKYeqMojg9ZJjSCF
OVEGnRtQBveH7Umj2BWeJ7J36Y/OAkmxANj9lx262F0AO1QJWIzoJL2L/cmYPpRgGoVEp0rXHnnP
Ab8CJUSh3kxVC3OcGNe3ue7pFLhlNDVv6LoZkp7URpqb+7Ap5srhfM8C2YZiVO9U4K5GRtY4iPgq
VuHAOZzvP6rDe9643OneYU97R9MDU6N2LVMwTWzwpZuuwRAdJ6ECD03j/GaDnAWQ7xYM5LYMDxPz
8X67ziCVhh/Dj2KPH3h2Jg9PaFUBdwI7uAznbWKmb3AQDxiPDZEIbnQoVcpD09o5DlJB4ZYn4+u3
2wIET10Zc+B29BztEUeiovcZmEXlIYmuI+SdPwGPFo6jh3sSotXfIJ0//hvZ5PyYwqSuFRMQun6m
dbqAJpaDI6h+EpOv+a0uuOBEhFUUm7qUyA4eDwB8BHqO/y7BZdt2EKC0JZ1dTa4lXVTlRBMCQtye
OJbpF7k9+Kf+Wy3ej6EejReOkjt3CVV2zQleh0AHJXXjnXAIsnocRF/PnI7vjJen84jJAA15lBx2
fEolO8vIr+KAsDUIuDxLLf1pxCwgKQBoKAl4j2hRkZVRpgNnj8sM1bckqhVuAwnz52V1spmLUwel
Q9ExhEpX5yZh95wo3FpdR81tRMYebA8SiBWMQn1F/Z7qoKMjNs51K+H6tZcArzIn2XqhMhsWwu8G
JG5ZUYwF2K0ykoUzzTExjXSRrI+QqWZ5BdxTjptmxT3Fcl+lYlxopNdCtQ/enmNiVHR3CD6Xq7R+
eB4/aUVKWVULy+6iegy0x/kUsbLnCHvH8c3A0s63fRBxZ2I53W2OrEDXuRa7FMgIT67SA/+Gr5tN
1zULjFCoz3g6lguqrWo+SYI4JszmVso1M5HB/19GYpSCNgozixma+c7KWepr+o9IIcYvtr0K4byf
Nvz6MUEkYrikEHfqmRp9QEfzcDauquRKCH+FaNdgYJPznD7+CZovcSKYp7VGuPozdfBGi9V/A3b8
YH5JrZWt2/XziuyWTVO/nvfRLcXztmQbvLzhmXOu6XvABi681ELciMOGMFkAP+cO81USLnnGqOrE
7NZaw8LiiizMW7WB+5omzRDZrb7yum35PiYJGvOwX/Oqd3fTxe4soVbhcdzhPmhpr8SJk+cE4roS
bVAD+LzuU+xTD6APA7bc+gMOHuqPVUw4uU2dbef/8sSuZu2XPfGYJIoreYuhoP043ieaMjZuq+1y
h0lhGw7eBZMd6/6u9GcLl0TTggENXvLrpu+Mt1q2RVy/uDi+lZqbbUg6kJD+NddygUcitV888MWp
T+ct6RvAuUT+mQu+BiVzQSMe96UQoXjD+g9joRk52eDf+dsmwkhFBqoALiBYgr/XewTt88UlALnB
T65w1T1FZvTbf47OrtLIgFo8zVP0qSbozGok53J9mE35y28VEIqKtpCHJpbQBtAA6Zfqo873dzOL
ADwKCA8HkMnyZ/Cqjvtia+TJ9m57ic108AtRhhKTZw8U9R7z8RWWT7TXWO0KWBdV7/QZ2wvrBp17
dNLw/SrG/jNCIKqxA1OHVsx3xM2xE+I4fS96GHl6NdX4y0of6WMvqj3ZHrLHbHrQQbO0GO5A1zER
JTyIjhtK7Pm0xWvwHA1a7+DVX+ILSbWbDMr0AXwznPF5tfivu3rHGo8tLO6DMP5vENBrOSuOuEx1
TCoFTFZckw2+slZpYFSUkPK5Hmzy2I6GLSSiqOte50zAksGXuBZKvcLVQe2/YSI0W8Ivqeqx9UF8
OGVUao9UgbxiXivHF8VqtGWiIuNhzUPm85QlZqxii8DUjEndEngY1SMB4Ii3JTPkufNhCuN/dPTg
TO6JnlqSYehJV3A2rtmcY4gCZxbwUHHPnxXNm1ao5w+abgKddX86ooW0WrODLS0jX16KMpAiJ95v
IqaoubpE3b/odpTA/zMZrWbDoYSXMq3GJYjHGJiplU/PGHv+en9OXS2TedOsU1PZn2+YzBY6HAjb
QVmj6JZFf72VE5sJymgmwtogc3AxchMt9ZYqTIiQAAkHBotWCpzHrJmuilP+Dq8IojADSOZhr13D
XhrJagBInIRmG4h6LUwSITJ+7+ra7Gtp+Z47rr2lm8RuVBD2JAPJ2YdboAHz8FFn17k29lHdf7bd
BQZlzRrfPRARiBEEqICvchfk88iMeLg35Uth8UCAzsXaX9tvAq58xTYwfaDKWJvqF0YCGzQCEHfR
Ry7tBbPKBPMsKJTIHEO6tdPoiJcrIjg0aUmFCjAZ+F4lLRTmADhC9RMbarcVWKkmxWI14PCYCKmD
WxF3GvCjyTc42uDBD3JZg0jbOVBKPx26CJ5HM2DsuunRbgm4KAXAlPB6h/WjDzElc4oVODmJhjVH
tvcQ5+hQ5nrXJIO2GvV4OHn9TFQrD/sT+KTy+4SD9de3uaIm7qK/DZea7kQd3Q8hVz1FNUMWy+b6
d11sm5HuL8dvutW2mp4xmdFp/0Xmarpkn+y6128lUoOCrgOPBr3+vYKKGI7Rhdn3FC8eTzj6PghS
GaGgw0vNiZrnPOCRa3yYRGVdh/trKQGbWsREYSvmitmnLVaDLKu9bC4trhDRUsAKGXLDO/yor0yR
Ss/N8lS2KCd55+zF6JsP3mPgxiauQb10a7LoamMInuZoExQ4a9s/zWPLyB0NSJLvYb8nYwV6lMfy
7OrBc4r4KLsRdNbbSYzBxIbwl7vl6a6d+cYd2eaLRBweJBCMhztu+rUFPIlijqLondsihdBEH+jj
ArX+/7Yn3vUYBYdwMsJx2mzJtZ/J4OPfPW6J1w1gWA8ovpZV5LVAZPh8tipfpSQS6SNxnXjGeS9H
q5OsRySkgTP8r4WplvBXT56TJx4/5CUexrEwrdoIOOUGzEhTUZJT0ytpkcSAhr/In6ixMSbYU5ox
yCRe7JTp7pcwTV0rsXmJFULFjpGTQP0lvda7nrDgOREZr1d33nxH6ye08QAgPYIZw3/IAHl/Itp2
eqo2OSOnK2kkgr+r/c13TOTLGxNO3Xedi+sKlFxOxGDvgjWIVFIEgeR3A+1zZht9NbjUAT7xm6C0
+m50+qE+Okczuy/UOkwQ6yXjlXEJZAE1S8kd1FKiTCGKYrCPi5L6v0Ib5XSWIQ2MdLTIjJfgXnor
ITI6244ns7ZuZjB2s7yF9RCKWkRvNLGgwYrght7hgqITYedBAl9aiYBJYePZdostC/RgtkYof3gp
332hAcyXiszunTX64MTaCOq2D+ewP25Yh21EFM4bEtUc0KwVSjMm1k6abIMBwFUBY52PfNdv4zPS
JtWFY+NJBP2ws12UI/HypqpMsNAMR7BCshPhsOfc8jsDExR4kFystQxxYp6jHa3tdaoCnSdfZvpi
4Qyn9Y3OCXN26hRKYXuRLnvwAhQkLKvbtbtTenoZk0sh0eEGgNSFk+DyYlhm9GnmwuWUThHfuX4Q
MDvH5nmw2yAMqgCAkPSKxh4VcNL4j/FIVvmtDwhk1iXMlCshro9uj5ZyyJSyvu0lB8O7YOS1TT7/
UXJCyE5j0irQ4W302tcGut3Me4mIhVUYlZXJGaVulEFksSj7h4wO2pCdM31EA7lJKN21fAhJtYM+
gfTIl98AhDYxDO/TlNaWvAdYtc+KTaN5ih8r/l33qNxnAwQywk3GniYgtg6T3ySbIYL6SW/ovgM1
qe8+99LuWZgqlAO3mbBgaIxn6gVX3PjCOKt71oQ/ZPHhw4n91kh+VP9lnC9p5Z3lnmaEE9HndGa6
YmWyrIXqjoilY0tule1DyMCHLyjz1woKgvISXXI6WQyyZW/oVbByArk4VbPcrpVgz5rbZTDewOng
4PNAIzURqVYd+urM2HNoku/IDn0UocaneA6YNJwkebl2rjaywGs62LYDiiIzS1/9myxe9fEn1b+Q
qDs0LqogiNTyCNV9oUJmUk56i/VhBcccq8juBD2lvAjkD6L7Fu4Hw8BBeTCD5va7maNU0N8mMUC8
SLyZflyRLpiBzhwpdnJtmVF7yN7TBh+rzaG0rpTkOvkAcNciCFOcTiiF9qVGTRoG4ArfgSO+pNYc
HgwmuRgPCqsXp9TBrndbF1YhgY7U9aDgwT5wPtICedzriZGWxgkpYCSY5oiHiGkf3r/n4eb1BP4B
ZbCDS3dfZ7x2RXJ0j1phlMmyPQzR7Of2uDxAwQSm2qGf/e0M2mnUDjmmEDXgO1JtY1afnMBbww0G
cn19fs8ogj6HNLgl2uq9P5mpk9bwPyEjvuPcF39RQ+pCrMVTxthLJyGcocndoWBrfIAp2hRwpCaK
jkwcIZH/AfxG7U0VffmrOQptFshw8m9nkS97wduc3XTzEfYSTktREZfH7OhVurMfi93VLptMC97C
2/PVDjiyyGfIBK/GJa6PuzPF57VNtj+v4RIUUID0vWPa+ZDyRUYSlW+rEfaM4RTW1tDOy5p2JRgg
lBouD57Fk2PaIkjdjgP5Yv/WAW0sw5Yyyc0X6MU22Y79tOgsUCFj28st+gyFkCM/VdcgL035I2cZ
Cp9F0kL1E0AvRrHZ4uK0dFyZOEzC04Qo4aeJXMpiui8qQ5lRuY+tV8YLMmIqp5jSWxFwwgbYvYTb
PXC2+LKGUIl7l0ecaCSsuAkV4viuHcINHHOQrNepDHBNkTHFoT+t7jPzTD6S9ns1pqdsWW7HEG3v
UFIRNBb1FI9GAPMUL/Ih3OojA9vToXOEn0097zKpmeBWWAqLDleskewFcgMnAuvC/ZbwOcXKXgaV
tiT3NTbMt5Vl4GXPVmQC465K0D1yfCVH+YUSqBwJ/aTQgbTOrkRGxhEGY96HACXuCGBvlkNiuzTc
yPohPyR9r6qn9fr/Re4IM104DtQDPsEzBt8dkonuO6sA8cLai/U/ZFDGTG+9kXpnE39H+LGI5fQq
MF9anM9fCiy252x8zb6F4+bGK8P0U4NEMGCasddPSPu8VTOUCceyuFgrS4gkBbEGSwHkfWkfEyQn
VfYGMpMS3fr8ov035+ujJfLQakOrtAgtxNbAzJRsW5r7SyALfcZ9LbUJTTD7WXyUecUEhZ4dbz/S
v8WJszj1BDkMonvlZlrZ+8MMmWsOiIi4aeUPd8mFEzWUWHelaBgRS6fWFqXGH8JOb4eb6dz7dTY8
skmH/PvZeQSSQnZDZXfKwKp4uZLr7oJSMtbK+1kVcjs0xmWS/tyLp1VoaoQwM1Lz4KNL+b1jG7oM
7BJyHX5iEr4l6ondHar7KLddXPGAYPCS5wQyR6CmMMs6wDztBVNl9nHPH4SxPs5yPgF8LrqK5JJg
mpVcaQoVEPk0d9suedk2MgZBbYvomf3br6IqQKOgEvlNS/ABynOCTpZKlWfatGiXWab+DQ1wmMBM
6CRuxmxeQfa1mYVi3iHyknMAytcZ79GRH9zli6IgWWio111OTjFd4d4/ci5kdgjF5cNDZvukD+ck
6DIGkkiKi2Tbc4ZXPMQghg6MFk/ub4uqWC02htEv/RSNC0HNLscZwdws8u3RFvD4yQqxsBle54LH
m3R0FaFILXqMfXgUAUFEtO01Xq6L7RE8aE+XO5TS3pJn9C/zzOVl5Lp/vel8jLYv5NtHNOxHJ+gm
582cDrOo0f4N/qinl89Qle1i4mwba2ZP5me8nWE9z+XgY/+c7t/RZkDSFWdKkFmJ0W9yb/yrFXyo
TbPOHbeS3Ujw5g1Unlwen8vKd70AM1KK5ZP3yxs4LiPVZLf4NLy63wq5PfXlBdO0m5sphwHE+9SF
KmuIreBdPJ+ZS+XfDmlBp5+3h8GRRIaHbx2OxqnqYLU3eMwTREZemhYBTZ1PhxHMUcvN+SB+VmEY
HZR0IpEOyMXQOmWHvAAr8+KmqT4gAMgHsFHo8a6f8lBiMZAKMkGkn+3v/B68ki0lXLc3u3kd+4Ft
BurO3BrXHQJhQ4vYdlZCoJdbqUT3SZm8lhb07NJZ95qxYOiHf39YTJYl8ZIgOeUfmTMvUj183hvU
d4qV0UTmQ/GkBYWvRYg0jz+sIp4qKTqHX2mUDBx9QnNkAQd54W3Q3oF9qn8Cs5w8Eftc07PtKlCL
tPYjMmKXjAnzjKmZaenOXmZ+YgFkK25EUBkRhE/iJFePG31laNEU03+rtIRSvXUHFEr9hkXwiEYp
bR9Gcp1E8aXIiwXl8t60zwSMxmyAc4MQ86cA0rpioPubXqnIjhHX8QJZH+8zjJ1F0bKVgzhjMy9l
xq1Fddvi8hhI2/cQBsjEaB/C6soI5xcliN/uCb6ajnEiBA+a3U/a41m6q/4PjetUD48cXpG66teF
go9xabs8jhlyJIIMC6IROD5ZGd5SayHeDYlGgRiX2eval2jXm57F6Q/cz65o18Mc8l1mG1i7C+Z+
EA2W2d1j4GM1GzaHTGWjvU1RvXQ9tI+rJHXRw/xQTpVEAuGgBKHNk3CEDDv2N0M/y19+ue2/S7xs
DpNROkR/ko69W+nUBMrgcIPqKneTWR7B+SLIao2aCzEU8xFFT25/cgPtfSeqjbkvRi+GL68gLKTo
9xzT56XG+1SJGOi2LYHiJtTlPcN+swKymYTbmxXOmWWgmTUtZgQe9chn92NnKWmTc8tdBFkNkIW/
Q9SuEVs0bH9VOzdKe1t4z/XjLDANPsB2EE8h5jSmyfnebDGVYQfQsGIGhgwCyyR/BzWeBobPya/V
+dviqGsyKepw6HdlAWqWjqZnbI75T55AblbD4yh2/4KzCCmlH8WwQtimogmfuQEW0RjGgCPrq30c
pMt6AURKAR6WWY8AOKn1pClprSQmQHvdz4oeSU2YxNuWppB5AnA/zRu00rxLNdoGVN7OkmPk8w0V
3VR+r9ghaKhAAkTyqFZIwQrkCz+0AKmKP1ZCN9UxoW4ewizXUFu4t5+/DAUqOddgM5yntlSao/B9
n40BNsLv+gmmxCvwB42K4bX/pPdvplogW/5BvLwes708/l0NwC/0x8HWMmnQl+jQG+nvmijfakbn
TkSY6juqDTS+h62GRXHFe/EzOVxFLBGq8giuXozgyKkHQopAKl6bNzoHa2BDj4WLJaCxut0XoigO
fdc6z+5E+OMdZL6lMBM3fsSx/hkapAJ4PpzLVpNUkSe18whEFeGIpCUrL2Vs3Opy9B7EO8K0kdZf
7PeIkvS7n0cL8ZWGiuyvoOTA0M+zlwFQSJO6QdU2JvapHLkYZHOljnl26mxLRUE/4YSZ5Qi7XN38
9mdHPlu8aAnWrVmxfeLnAVT8BynGU8AzLnrc9dOrrjbNaH2tiisZiGJLHDQxiJLYw0K6Z7EzJJL9
azXLaxCMbVAC6qS4jlQRbaU5dMeBhdtP8db0rRnempkcYvSaLrImiqGnH2KFi9Pfn0w1lC3wWTct
J9KmkZPPMz8MWVRqzYQSCVO77CpQgJvfIWMCPRLpaseHJvnMXHHNjkUTaPYsVgKJ+P+O/5fjd8f+
jtYLVL27vGJqRbzgkRKp41Qq65Fpds9g3LX3SKfQFeWSXpmqmrlfiJIJPC+grjOkDjGurmm+rAbd
yPhJodlY9iro09tMIHSk16zdAuCFsRDNYOO21fsJBV7jC4pOgncnBU+vPAHAQGYZxUQXdFbPT+lS
kRfeNFyHMxoJQc2accrGDE1gADUwXti4jNH3iqWyY5mmwyXM/AUPN9SAhtvtkwnzuWkYLlLGAG0d
luxbEFg2wi1eSqRFxJM/V2IpvkaAlf/2OjRY7XQV1q/sFLbS7uTv1G3VbE5jxxfG8ChlfS5O8ubH
gfKWEN7K2ErTEaOW1qdwFnL9iuMZ6M2qLCxaSFDg6Bz+lB70hCo3kPwnxkHIpgczsKgkj4eCjlrc
vH0Ah2ThWdlF8wQ9UJJKJCQLrm/Uen6ueYqLsm0XW/34uAU9n+ZqPmMnDRQMRbaXTOZsbBkYs58R
118kB9pNRuxMI21GKzydHYEgeFbsckNgMFQLLlpRfhaKp65t/G/uYgUI+xwqNeNHt/GjfQvPTe+B
REbxucVPM205wAOdj+/oWZ0tQEeKsNt+uY0kuXXA67weowhn6mjkJ9M14jrDQTKxB2j7xbosk/Ti
GQzIaI2CQoVU8Yf4CuHeBdZfwd6DR6RilbCey1su2Tk78YAgD5NbXSCreomVLon7hBd48FiNMR3v
oXpTvlWCbzGpupdEvMBlws7h6D4UtfiyA6m+YRJE9sPnCUmgPVR3qLOBuOzlAglPZRegQaL/7CwW
Vf+vfF/X8+JrQ1ucRtgRrOtMALoiYNoBf5uj5t5K0UGr0IvlZno6b+judXeTBO8OF9NWUgnkDO3J
8ydGsJ5lvxn4V5nO/8/Ox27DgO6tlIMFcxLBZe4+xtk4Fbwo64TYsZkU6S+YnFbC3E0IDAvJZWH/
os8ZzTNetfj0nOrDX6bNx1qEhiM5zHkJYsYcJJvA8kqW5AC8Jym/P5OmvchBSz9x6wuj28XQub5m
KvCHLtfKHfGRw5MGSzh28btbOwON9mAzLfb5Us5Aub+SgD4sFoSnJznIG9ZB56zQm78n16FTAX7c
tXIVOAnJvkdAFl0zc4xWs7HVLCVDAlo/ndkhXN4TSfhHC05qRV6d1hzS7tqH2wNMn1mNwh5e5yA0
3y1YHj6voPr0A7XWBxsq3RXyC0JLeemlJLc3lDbSO0NNs1dUhYRlcxH7YJaiOxhLScqhZmBEFcUj
0hL7vc1J3Wf+yIb6lf0O05OqESBezoevuflGkuxEuE9TPW7iuoNQktOc4soD5vU9nBhabi7ddvg/
u+vZ1hG5LpO4VBoXFtmN++qHhzSNDOWDvvUkRPz2wWdCXihvSokhlGVGwETNn/KzanqBeIi9JrmD
lf8bDlns0Gcr4YyryWPM4+eQvM4sVTesW+zGSH9qeit/lykD86EYmzGs/b6nVUD+xY/D16vQVgYl
1JBRSh7cCh3ky3DwAa/dCUhiFntf/FFw9dRLgGPAr5BI3APpPyMvf0t3SoimQF9Fhu1YHc8MfhBC
gH0F0XHNJiOzqA2fFRK6tVYzX1pAV4scaKLNxQaAdBVh/nGGskwlJAdf2qO22MALuaKQjKA7Z8/u
G3wknODwilqy4Ww2NS0hKeaym338J2AFaqdzTocNMAYmlPjNH9dH4r6bf8m9pDIgzO8peVX6nAW6
eNpTALMqRk+/3SfCcN7VtQLYOdCYljqgPFn48jF14nQ3PiBNtnSPH/8QiCxDFZ93JWzg/OW05hT5
+BQxgw1S+cj1T0P7IEXnfxuQQ5S9yAMvmTdKhPAJ1jpNdKbbEcJ1FTR6PetFRTJ/7Y9mHjGHM/p2
ZqNHkJgsefrYaOfuvWeSesDQDhCYnaA9jOH4iy8RNDRd3hjLruAybl8Lpzt/DTGb0LMILteavLhV
AqTP6VoM1SGTlfuvO9ZIsr+YpBxnJltJGndVNyLCVva8+pTFGEUA+E3BY+WqWT6hd/SCds1wk4YY
m9V7mwQblRxlB7zB6gAxqzLybHwJnHnYcT55pGWsEoQnP4Zg2fZjZHa8lfgukpEWG5vr5Vn8MTmh
9+WDS3OswAU/J9y1iKW/4tMmKoRFkTatld+xSVA5QkHk5VkAhZzJIICB+OoGiSEqlyF6kls4x8J5
9HaZtEoQWsHhdwb6tAt0DHlQ284gjlFRGh8U7oU4sfXSazfDZ+2SBcB6pddAiNdGD38bILXXGC9E
GJE5V5kU5QBphjlwtKJEOBTvwNiK9PNNgDmlIELOgPqBKNdde5NOlesbXH+lQ1mmI+GcmGSg5AB9
p72UiKv4HgL5b3exGq3Ghzn7vCp/slX9Q4g0mMaogf2bxWOjevmaOFxcwrCCFbwI/ceb9OeDrmpA
cLnpzVeuGzs21pJuYB09I51vCzBK/Vp7+zEWR0Z4WN5h7fE4efFxHAOTWzJ8RNnOAqabBTnGRy1P
7Otv11MUrCI6DbANcM620skE9oUxaoRyilRvRj8nRyq3zqmmYowN3GxdnRAc/9LtqTQrb5+YJBUL
rtVgvjoYtR0Q+c4LTi8/RN22hqXnp6irN/DcbtQ0Rs5XF+wWBVURPJDtiPzo/XEHC0VANO9xcNCt
XszfQX/fblGkkRChWJiAmAZn+k+TSTSJtP7Yvc6QFQs/8LHZ8PcVnBM8y/7rtvH+klRZPtKEHRk9
xi0qGNiLnBb073gHfIYrk3XQeU2DebggisnAXTNgHHBjQt9bst0qfiXt8xuvQhLxJZdAhR2O/fr5
Q5de7nPD05xxt4eIoiyQvhseklylS/Xg+XZS38KbadM8PPQgGzIEthGl1j4y/YfxZTavNdCE1VxG
fmjE/Q938n5D/oCZYi2vpJd8sgby4GODnRRNsh+XTjXM3XUfFsl7lYfhPXGXUeJS/va7D5X6bnul
NYGdoxIxUcaE6jdf2fPbXP0CJ2pi16Jm/NHieRt/zHWRW45GNhPFml8AvoCjeQV+lb22UMe3o2Lz
MBx+oDTufz8sKHKCE7b366OvZSlx1aLjNMJt6oYgjevvqe670Xqb62MN5xAfTaDXDnMPa2Dht5px
e7Zk5U4IYVCPTx4kZcdZ1XR/Mn3zETIV5K3cAxA3+q/+PKpw2pecRVQmDsaDAFBkznZSWKblRM6k
zv85jye/SNacPhoa3LI1jgQrZY8JGabwrk8apsc4z57WujJSpzxcYKmWlvOS9/XnMAiwE2C5pHk8
SWztta7YcZgelXNyDudu49HjB2y1c5YKqfi60StJGPpMkY5KA1NBNrJ/iVWArjUmI3IbWUsbM9Mk
jjsXhyrAIu6U6osIGijrQVhBZet32+jBMlOcJvRQBIRlO8q6PW7bADmXvTlD8SFa3ksCq6OYw6gT
1nExkLtPSIGkfkIS7c+33gUWcukP+JOorL3nWhqnneUSgEb/rtv01sZvE7P17duJ53qHZeAY3UEd
mZ7zDrCfxtGWYvL5gbsy6lyCuo28TY5IT3dY266QFysK9XLzDnbysuaeo5EkB3hnLQVE8rWF6LSO
5uC4bgoRdKnIv56SMhS8jJo3snf1QcuR7Yz80KEsK7EF9hTGYYEaZcv/5I/eoCHnxHLuwlZYx930
EF7Okt8TsPuSR1xk1ijw3up7yVrLJSFqsLrHWGpts1n0AHPCHZEsqYx3M6npI4lx+Gn8vuYhA6Tk
A7to4SYWHDix7uKbWiBWD7FO/NkGOEC/6OCxmF15Tv10ulym4z9u5jC+KzLogQeuszDa3dNxoNyN
rOOlc0xAtwY8BktWzezeAT5G6ZDR25FyitFSe0AdWqjmfqHHCrSj/4RtnepJti9RIH3ruliZ71jQ
lAvFMg3PVFr/hRdcf17aqE/8bxpFB6Ws1p2xINdAKt/XpDhxfFnra7Y/ZhLftXetWQyQy2oXxAvu
u2FSqoLX9nkRV+iYyGj1yRlMPTyIbU2hOnyr3NPPl5KIfhcZbg9slLiE5OD6J+QOB6I72M7Dz8yN
1aFFS91aawxI6gc/+L4aLJ17LUfOyhWeJptZZbuUloKC8L+MD3SPox5NUUjYXDpbZnps8Zy8FNSE
dSj/ouN2cEKVw4B+ey/UiwIAZRfCbXRy+dHg63JK2O5rGx/PFdU70q+PmCxuHXbuK7GU85ahNkOn
KyJ/lCKdPfqJSGgUkEEvCIJfI5ESe6Az9cEQKjJmkb79ptB2mSHQwFzPa9hitlmxbULmAA61MPBd
22lpjlvPGJs+tjxVymFkx3aArijP4BVQfgEAd0Ck+JK+iG7+eLyG+ATsQ8lW00ssty6K7Hg7ATMa
1RFTC22t+7Krzdw36qmWCukEzql44dpkgCH3mAdQ/N+jrLwJP/iQO1OhejSdWg4H8Flik9pc0vsN
LMjRGehr/QevYY9GURjdqTehc3qZfWd/DfJcLrjGMWJV0S7nTfE+Bpcw6GLn6urJQt+ipgf9OfVY
8UDz+AjVbVARzb/q3YY21Fz4mVcJeqtA7AMfUl2Kj/8nndSQ/e37K9/DUCMTXEJyHE9X+Vc2249z
l5dn1ZD6G8Puc1BQnxjQwbvY3SFBkzQGmhgZLHfRTm4yt8JDjG3CdnHarl7Rrt5+2MhifVi7cL6A
gk/yhPsJ0nJK6sJLiCAsGxWqZ0yxiTLY92ElUl2AZXQnUBrxNtmc3BiJItylTbOJUCqGJCppmuuE
XItQ2GuDl+YWv3xrCCfskydac57dNFh6yMMJdNjw4d30NWB8jvII40TYXzpcT4Ekgxw3alsEoWKv
d5q6I4DVCQpkBuqdlfyp7LaOqegp1TTlwk/xzQPYoseleB+5aJDwufnMBrPOLZxhOSo655s0419U
e3p73DyuwPJGp+WyuubXyso5KMAHgGlGA1OZHG0Hw2FI4iJBBDq+KIsbYVe+DB3czZRMqxbcuhL8
6qRvwX8U8OewhY1Yi4EU26jOhV1WJuomM4nxHS/ZPdwKrNzwjpEFFUQSrgcDXFlw5kFL9hoJhDtb
DXDfKapgRUoSX7SHvk5KymY2pB3fQPUUjwRFfDv2L2S+tMGj1DmP7xVECw0Zzr01IFu8PtoGV0Na
MEskVBYoEFv5YJnk05v1/MLxWOlzjSvBlBH1Vbfc+vlA9zfPHoo1gXIpQaxkO6JQSMM/kYeLWqrh
aXWZKmLtk0LvlvguBshqXSaUaNiZeSCLitAvyv2NB+BakI28oiVotGNHOPSlZRXWMGMCGVX0t/Q9
sbektgfOgT6VEWi3zyjiDhbjya5PRw3TLHCcxVmd6zmDgb+4cTZy71nUecKKCfpxHJ0yCOfwXN3R
eE8ICmBUZmzicOuKMsMAtRmrhUtRoe16ZsBKCc8slCd7qyoBfLl33mrEIP3XedzpwrWOayvT5Pz4
dxPP50Fqr28Ww+pQmQdmqWqZMmpqDKEqSt9FwQQQGxAdGV5eISxVCNAEPrPmC5866OGK3BnWln4a
98iqq8gXyKrCnueZnjyv5OIu4HV6EjoZLHlk4ulj0oRaALQMZ7Gbmo04xVNqJucRFrup3qjTFGdb
ye8yG6wtccvDLPXjVRTc0ociv0NfJ11BBbnrVYtfYzW5EMYLKy56SN67YDSJcI5XYpHM7826Gcu0
xTA9gVH6J1bWYcJDVfbBlyXvDeKbdqPogrp5c96TDs2BtpWPrpY9tsZmTSttKU/9rZx9irP+o3bo
rBzF3iCbaLXeY/gM/Z1L9O6ZHfXKWTaZYBlZof2T3xkLcvvX+kmR6MrCmk2oimNkTtLOZz5af6j2
bFH8MXmh2CZk/JgC8zUA3ji86Lffy1oN4UFfdAWwx/KCLxugC7SyQeqFa40eVaVFO7GHgrhX0KH6
Obes8j3we1QdetI+VlGhNCswNCKpqyCoxNH+LoedMcFgZ8wStZQzzjqVAsHrVLvPEHWdWWnlnXZ5
CHVhXgxm8spuVk5AHD1WaBJbXkPfjmlESkowHxoDZWofBGFSnyQh+topzvAuPHwT/Ed6yYV9hqTZ
TR6o5jqvW85C7eVh+CdcBNFVzfVmw5eiCqzenfhgdx6p8PqzzUUyJV7AslMMp7Mp0BR8B4j4pwWg
oZEK6tch3QBhsvCX+w59w6kJEN7L85MYl3PlyybuJ8OmygoQBEPEfSVLW+CMBW9kbaprWIHXFPS3
oO9oNyltWRxfNPCiRvDy0wnPVjq7fzYUxygAkvbVzNlD9JPKeImq+kKNvccS9oT0Rno9GMO5ba8f
9OZAHlZzxXXNISzrG9soxrm8fs+EyMUhCKY8YI7gxOouFbPeTpvQ00YecqCJFMKyIwU/XklASAeu
NZe4DuXg4PwfRffkbQJvYNUvcThwaTBOh4o7DLJSPG1UA414I9eX/QY4KdR3HxA05O3FrI3k/ozT
joGZByZqqz4HsovQsWLqnBJi725C0c4mcmbNmEnh7mLqZBH8IfoMwpzMMtNxQXtpYp2RJCSC51N9
tqnsjQU6K1JplXnFJVSx9EjHu1jnu8t9DBbDLD10ApFF8uZpgV6qFr4dLbPMCeKbrtigMquupk6C
+PXwwPB2AhHuFd2yodwgFisKIlQZkAHl+PodiByv+/tkgoDl6gl0bfsC5T2ou3R/2BFjEIEePuyQ
rkFOZEdkRItrIoOfnBJJr2Z/rDfkCTLAnD2HQn/dQ+TBrSA3K9kvJrZRMc30XfQTvAWSo7YEyDbd
Gdqtgh3vlw6DCnI8RIUNPXFw+wyRJcih7YzbVoWbsNYlbrWSWihM5CxDU840vUG3Vf07QXpCLa28
+eJfz+IzRcgzk1Or81X1l6Ww16GRIhsM0hed2bfV3rQ23MMvXutbH5ZmqtrbpOHsxIRFXGuzTw5v
LEEcxmI0Uo9Q1r0X4yoUE7YGMiS4SDWimcLhiZYfN3IOWv6o96eyAeFedFq3ZaaOF8amKuUEHRlE
6qv9Uyjqpc/61S9qfsR3jnqeI5MajKWNNdD/5lKT2JB4DZzbcFDbhkzmQ89u0u/+I/xLeWQpRlb7
ejk34Aw84pJsQdhYURxFr/kWRzFBAMl7sQe1aqdiY6y0IwJBJIp1h3sW4wNhR+Yc+UGhuamiFrpJ
24A3vY2n+d3pCC7ImGfoWI6DIS+MJ2o2UPP/1VsyhgW4avMGp67mM8ugeA5/0b8h+sUug7RrkxNN
Ef1GS92nR/NKys6kfLLE0b1tk52NPQ113BJ8Y+TBQWZbanZOfaCN8XsekcW+W63rHGP9cRQzgRp7
RIaeWG2T1ltUR0DNZMVet/mODLp9OZ8yZ7Wsl+zPaak0p3nR3iG+5xnb4lvW2sygAfsM/O3gi5Tx
KFMFSCjfB/PmHrXQxI33BIN0iP8P14m3bPqqpdwZdrCKhcMAOfCzqSk3eOW/gD3Tse4VmFgyKjYW
/vuxH6M5qrHz41KZgbVfdESj+LgQh7zGBQDvz/ewYUR4nF8qMvVzXHnDrJh70NIppV5w0xfjEqzx
CThCCTp84f3PScN4sbk68BBddqZlC/8k4H3VznqmoBFGwrN5pIFyq5fXtxC1LnIGzbefpmLZe9Fd
JKOwLZ7KnW/GDCRt4LnBZr/W1Mn76sVG042zaLD9DHsSKziZsXWzTlcnwmn/cOFbMlZLSNYh0Vnz
bVQqwLTuKwFCyS7785tijgc2SYfSQxhDw9IBYFO2ohXd2/XNXdtZXoCcszdTgg5jrTDOPnNJaLpJ
gXGWFK20mgU4wtlQbJoI496ENai8x/NoMKJRf12s0dJZ95oFRlYFHdARr62feYspXdOGuFwAG4k9
MkLYKU1U+y4OmuyakFjiFX6tgVvmyCitp22z1csSVyklBNio8BnIIMLnifLd4enWYLAsUo4L1flF
oeybl0k5qMEujnsjrWHnQ0G7+MWctsPwDczNGo4uxuMgXtnu+x8is2E8WPoRiKtb5mTTurdfhAQy
OUCWzgZd3VMdXFMAfAeKPuXHtg2fIBBarSOQ8wk2HUfRz8KIcEwgqrVuKOMcIZkuVsNIB3JrN5d3
GaYiDcK14oq34gTZN25xBBDJKTbTYP03KaqE1mdpdLlSDSN8nJn0bcuLYPTnecrECHoN/QwlLSO/
VrNf7TfkP40Y6CPZiJFYSZs9Cti1sbACBANR1bNJhuKPVpVkEDpmnTroUZTuwlhhBP5ObXIUp+s3
ExaxViyvHcs+VEI1DBucApq04IKMSAwPKzH4qWBWWfcH9iH3pDnn8GysAlOthZoBenOUCzz9IoPG
wCSz1FGsZGNsuslLaExi4wVndSo7EMwzFMa6UXhdQkDCf+lgjpcqGVOXjPT+Cq5NAIyFCN0Bx0+u
nCacd+VkWxuAOk7IViME52yGJl5i8wfNMuziXnZI2e+TJtwUfxNhdtJb3xV9iC2HXJPO2TD4no+r
0AtAxky/TGTLJB2F6I7imbUwsbO/vYdL3hPcktcou3Vh1HyOWDBmKWYan6svtr0ncBKCwVOVpRar
4TXclL7Ew4G0q+jUcSNuM26Qxct3AHmhYxj4mrVRVYhnt9KTRPDwX0vuA0stObWyu6CQtEsYm7LH
O/rjCYRT+FUW5uuXpAB1NT10JI/ziINdiEto+We3XbIGTEwHUa8MZeJVS+qbpukVB291xO7M9Wzu
+88Q4u98wnN3WLM27aGYqLagnXxF3atylM6OEYenroe6uiy0llQu8EL124AvY5/zUn1WtrIyjLU5
lzFjPQ2pAt/99lxAEtBrryeTVbxQu1bocb9RWjxiKIZjyk6uZtIKGlbsxeR+b1wtsWtBH++WNZoI
nEF555+C6rrK6pdRVgF0iA3APJOEmren3F6VRGDMka47KofgwwAtBxEW8wpIlJFOPOfTCnZNUFqC
3ONCQZYa8dSOI7c1GGQJvyuyjkjhu/uGIUtCiEl1lOAykHY3XlXNdbN11OfLRRXB/IcYsgiI1a0V
VxqY7/PLp1XD7nEcPS7Xtre2tbrmq4tzHfdfSaqdDWsjQovvLcbqOa88dp6YUHm3MEm2B+p8bmLO
GsegifFZ/iYP5AqvouC4bGnVlt5VNb4kQYfn0Y6li7WcLsJHFPmnv77s8zHPy5JEyYLQDjPag1eA
2Ee/pULvcj7KlbnklDG4Cz7KeZR9ik9KpDNBqN/KIBcIFCP9l1Ox9bcEZMvAPemhSM6bSI2n20/3
k4q51SvK3JXK6cjZ80ea3E7XgKUQPvgUSKB1OshUEAS4yQqsiZjfmm29/u8hYrzIWWqbtEykj3ox
IxG0hNo9kF4OrJD7PiALswxeapCGHe2M+oFikACZOkC6roiV3Ec223tJdU0pCUBEFdIIhUFZ0XSC
svNC7IOIcsHq4EY+OBF2mZvzU2g/vzFeoJIvLPMBN1iwzTe6ealr0/RJaZQBjlEsD5SYYJEVhWUQ
c88Y1WlSiVS/0B0qaK3dIvhYTCCkQO4iBfRnt7YTLrNBJILj/ZeayobPHOw3t1NMJPHI49VDMFIl
rYbbIFKebD9INeXHI5TZ6A0MeVMUZ+ZqnmU7/cFUggxMKzfRVxYZYnLj6LKExXVw9u0BtnoEPi2f
ivsVeDZy+dBgTFaYhewOMM8TYbB44j50zMh5C/uICbZbqVsswkrOFnkRDalHkihnR8lOHWiarwrA
mN/5wbyNLD/alxImSlpsaK/ylu8vJgIJX7ZPagcxmZWh2Lt+qLkpq4iqHg8NDrKCOh2In6NfWqgK
yEr73AFjpTLBls5ExitfArC/4W43YVXehXcFXLCMeQXKH+ZX510ep1YxqLXp8mjGTLxULx56QFqW
U7/HPGtUUOXbrpBWQVR7z37vJkHrsygq97sUG5UezDz7vq1ot/zkyZApWkUYL7ZapJNlY3kqFoRJ
WB7JXWw5PiyWP/9gn4jzoPF0hgmpC+qKyNlRPHw4PE08vBgFuJMnMqRPn9P7A6tlwmom6kgjPN5L
qGwN2FhUTquBGku6XhYJSJ2xbIOnXBQ02rG0Turpis+zpXXuKH6ZvfJENsF8AvK/rF3Xk8RhkHLz
7Tzjkz4lkkF3ELneLY+LZN5KRfCGdqAenH4BXask/AnyKcytf6eshxrTpRVg8MBSAc6e/tQzlaB5
CC0MtbASxFkZm+HzXn1yrIU+5bbXbNaIXhSBbHqQn/lNfaGoYtlX4rK2HdAuAo2QMFtjp0vWBKQu
IF8bXwgvnX4t4epdS+d8YzqrFyPYra4fSON2itAVyTpoXbpslfMg8RVVXpAODYLnsVGDhQQHQr5s
bjVDy8c8RFKYUxXYwdDWriSv8sEtbwZsRHcUpJb/nJKE5R0QiVK5sXFxW9cjaH/3P2Rjev+V3/k1
Dfpf7c6plGBrkZ733crXmFsr0QeJcLyuS7P8UYSDT9TfGDS0pG6Ui9J182UbuQT4zOhsFpD9u3jg
4rPqNAL5wgcubLrBBaXNlgrmpPP8/yh01zLIzf73oc56VHUflKB+CeweJ3T0XcEOAZeEduh3uJ4C
72DbHqhtLBguUQJttJpXnkLKaQp1bI3/j29zMHIoPZ/Ct7unmtAEcpycOXOElceRJr4jHfjqkKXi
zqn1NPupFHPA3tuHColOR5yVzYOA4JkWdYd6kynImAJVVjwZ6QWUtjVyTWXYnOJqGUrHqp6cB9wB
hWRNW2dKFeeBV7OYIpIaH/yFNNSHr+eQneWP0VzZxW2wlnHXes+od/QmwdaK05Hvj6L+GY/UjtF0
lk+xg0liyb7Ra59E5PoIhCa6lqxcntGvLNzVBmhFGJhUAbm/aaqkQf6X5DbSRV7RFxnMSD2O/4w5
jkvZy0UUJ37sfEi1by6m7N0oRb8sJlTqkaMVk8iIIDlgmxxSHr5j0b4Kqk9ngMWB62dDRU9dZF3+
HagSeM7IZXix4r4QEUilomg3up2Sv3mAAoZp9xiuysIycVy4Zg10XKTf0YoHh/G5SwIzBtDBglnV
lijE2nl/kTZJ9Ym+yy7jAyaK8+jPgK2VNURC4CNg1efLKSqo43A7IAlXNqzR5bfophjqVAxIfA7Y
YrAcsXbMUvw+Tzl4RssYwy028G49YbwimTbwI77uQBA8K6Wue7izFIoN1gjGitQijRXZY6NOdzCd
5CwfzCdA2FIHwlKPo1xcRnHGMV//8az2oj4YOs3Z2gZEewcGPEBw9vYqjG+GJmUvU+kM+GpyUgFP
JvAGgD0ccA+mol18dJfgxvrYLzt3WpYHfp3ConBADd26BU3H09XZfiVoqWwk1AhUvXnbsVc4P82O
Y+98legSwiI4pDBgPkwr6j6Alcv64NJmUWTzvHG7sKXfAV0UuzfQ/xDkIkUQPUc+LefJJEdykBhR
Y5pfazl9TshqB6dBic8EqPL2fSj4msXgB7d4BvUD2rJIPBIyTYMbGxg+4RVvGOITSnd3H7i4qV6F
luYR4vV6GDX/dVWmwgV2lgep13hBbPALXfo2nSoB7HhrecqEzbUzS0QCiUxQbUqlsDtAcbOqDYk/
nQHaGA61eG/eMZUa703g/DuwTz/AaRnoxD/Whbd9y5NG/s3l71JDSRfXewTMnovO8c4h1Ahm1UVo
SgmKn3mARCv76Imz4e6meQdZO7dbjpPHa17M0+BJ8sKySipdZyDMd/P4Z0vHLw+d8j+/ST+r2MC3
Io7VZxIfP3I6QXQIYq5d7TE9gl+PdLT6VpfKLpgu15E+uE7mDvO7GCXbBVTEnNEc2tv7xBL9/1Q2
GBpm4ALvejdj928yYD73+ZX43NtL6zLdmeVOTLyEwcgHCHOX2dJS+BMGYLyViinz2Ek/TG2MV+h9
iVimyef0XwooOI1daXMmuXzCr97JIccFz1NFvakHsYtNXwNzrv2jKL8K6jjTTi91f+//3EJFQ0zC
2tZAoOVneTOkuy0iu7yKFq8cEzj+/MXVh4J/PX7yTWjPn6DfnWwmcFA7/4fpItQQy7+Eti1tScx/
+UCHVtRIgto0QpzQh29jlbx2V0DTlPpARyyCtJepGQRF58T80FwGii1x37WsMYc5Yq/ckJEugGBi
FLniurJovLXmfNQZXamXpeMAc19RdqbuNaQ2V8kbJZLRx3Oy4PgEll1WECbvodBn9Xdmgi59l6Zk
hoEQhLl6m5F9cxsmn/ZXrhXbURj/qD7AgGWPTffF26XtwTr+MOaep2JycEMMDhnEyv8WLYKHfHIV
TqLbU5V7MOsElVNISajAB9aCkebHqQcP+92zETWamAgeneNtAL2DSdZDq1K83UHvIn4N2IJLotei
8NOaMtJ8EVfimAFEKYiXzlPo5JvTt4AfCgo8gMnq5vyF0wFQ4LpieFq6CcLTOhhNBABFxg0jQL9e
l00FlUiIl1Mh5ZFoCfvzM06HgBvRKxm2zQ+r8Q8W+YMGBb1XDHhBhLYNFEpJYQThlcOWhWrCDorP
sP+7/2lRu4Z8J/yTv+Op9u38KjBdS2x7Nbg0RSya+gXymtq3LI4WYUUeqhQxUn0gmb2WooocuEDl
Uwap4LzYll6ZRHliNrYfDS7J06ZDtT0pLUl8HMdMprm7Wav8AeUp1PjI94gVCl/cu/p9yMpUzg2h
wX0vhiSK+6ZsNNcWvm5Rm/sQ9feW1n9Bf91gG9z0lk8Xjkw58EcZERE9CFG+wFMaaEASPcHpGxlY
SPL2x1IOOa2t2xLbDXhp6cBlCuV8sRz3zZcgbp6qToVmF5bDGmuRvYfTrEPaaNRQ+gqDT+DOmkAq
hkiJaEPh63XEjyZgusME3LzVKNY+RqVUUCDzH41w8heAaAbGb4Z+0No8hZnbJRDJSE54h3sJYLLj
599ech9/tAqTP6efmbyLzUNgtfTju4oLJrK2gwqs56AwUtwNd83ABLog34lehrHrDGU31aNWqepa
S/LcfcYKVyoABHiN3ProqFOOBRd8jqHc6PYPS+YE4N88krkUFwxian9YWD6mqYw8hO724HryNVtX
U8RX68THdZWb6YnSEmU62o8JhJLhQFdcTg2IiACMu+5nS2go2P2UehfK4ng3Uy+AFlxUgt1Dar91
IO2qLnUVeraStgWVNoM9mhDq2dFV51qXSTAzdAikCAJ2BEMPFr4yjUwbNBGGcnlh7IhhV4sIab1U
Kj/D0hqXUG2y0kQY0hjpuhJ6Zvw71I8SYgaWFGeGSAY9zouBNP9FEBiM6Bb7R1N8jT1s3XJBj9+/
ctYtvSDis1sPT9+8ZwMaFl19kOpZ/SuxlfXNqIP5vT6TZ1oT0IqxeG+mT35JV/ufq4rX8LgOuGJ0
27ulHpBPeDRL4DK1c3UA3/XOEkt7y/knVExuPqH691Avdx2caVbqswJancOyEj56jUAqKZYBWqNA
DDa6jJgOOzWcpaBqInH45t6E7ex5a6uJJrT649Ov0yYbxpmVD/8eqayUjOvJy0TaOZZ8Og+lfMku
yHJPVSVwxGRepGuC/gRkSBfHKo11QMyX8mlf7cJ467nQ2m4q8p0jKbCJyhgaseqjrmNC0qdpcweo
LGD1rPrpVrwzTzc+sOWmlVtQLI9K2D+Fc3smuQz3vpCov6nGDzoHg4Dblgw2SWg5FSWsv1tNgYKb
8ly1SZ5slk1N+VjMxfcLZyO/rKFgR3/ceD/GximNJp7HGv/4IkTZ7LoNOVnOx/ZLZqH619Ip20s1
i0GjMetxWMuqxvXVFvY2ErmYG0mw1UuHdqZh5dgcxJ+6EI4B8uwWJoWwuwsmS141SqJw0q1fbICS
bmKxrFm83dcCP6Anxsu6mhIkYuS4NHvMN3qeJ70ChmR7hwVd+lLmpSD/iD4URsPrLVfy8ts0YuBf
uxa2u18urLLh0xQjix5oZmOm2t0xY+syPFa6TuwEO+UPTrU6KsN1+I7Eo2Oo7vOTzYDN0m7UCLWK
AO2lV9cNh+9yhLkJ77lhVJtLBLkmHmp6rn+gkm2F7IEc73WdAz09T17fLExQGcINT/ATJ5urqi8S
CXKeHL3Y8T813md24kh5j7CtKYCvMCZwWYHSsjeF4mqNPEy9B22aasAL2azJT6q6bZzyUDSkVVvM
BnZRihum1aX6KuXNhJd7QNwGnxvV17dkmQihCgnN5nvUu/tIFvDEx75Qjxu1ErTgZzh4MI7sWqgV
LE8yR2igwvJw7L97hH0K9LlnoEc4US6jV7op6T4HqjPbF0EayFvavnVTxRVciFmVKOhtdBZlSjke
wFudvHVicADY/U5s+bi90SzelmTSv327JzQwKsyiE1Wq/lCYxFWNgyDHgbZEucj5AIHqijidns1E
4L5PhmPQ9fUk5PF8O02F3xZWPd6LGkZ0C8OyXx2kcaAdrHqhLgPoha2+FRmbcMPvwgZErkQQk/75
r6I0rn8A8gMSKTnUXGi9D+WT+/moftGV3PuNm0wdzTNGkQmlR5B5+IKgTV5tKXtmiotZ1X7WzeCG
bR9sML/8fScsl+DeppSamqJ9aVeE4IB6tN2yerrv0hm8cmGAhVWBpC31Uw0R2+cnSJZuoeuPNjhH
bUL3aBSI6Yjp9WHCSaulCQJNL6ftVcq7enmUBpk4yXnoET8bBWHDXOp6xByAtHf9wNMOR/FK2A1a
ZYi47+XQInD2xbzQXzzRqGKq1XzQbGKn+pogRWmSD6pX4K4jVuZ5L/IiMJxUXK82VkSh0zUS1Y2K
+903e5qO7w8Wglsh7uX2s6faVOe44NGDQqFy9Tr+9xw1rTJ1CMmLtbRIIpaqGjk8lWmfNKmAaYcu
IUGBA2pHyiMnlpGYKkkcIZBo3qqq/LgPONxajlgdy+wkFiEk6NrS/bonb8BIA2NHBDR9340Bskzz
LHsURNXva9v2s7UFjG0kuc9UqJwAZPVfS1lTFJl+SAVLqih7K+7xgWND9TzSVHnW0O6+fu+8UAKp
OWwvlGzzrjND//XWkUmUgR9Oqm4cxHZwYXZH32JVozvt4OEzoB8o6aQ7SDBNHwgSPQVxkh8W+6Ho
4HAWBqNLKNdl7gCRVl5cPsyL5E3wupdVZryKN5dYeWgiCotThyri41xY7uezj0UUOV7MrZcVn0bp
uzpC7KKjqJfJITx19RRppMtdvUt8IX6Te4vwKbh2GUO3OGAxQ8nEfziGUgALRPU5gKmoQssKqDLE
eIEmjkGKd7xBYVsvqqAJx6BYeOHLRF3YtOGkJZvrVhka8ZDvJBQxG8zVv0dnsFkWdKgYgL7tsnTl
kkAvoGJES2Z4lpC+FtEA/vERN/N8r5EWW3vx5UTIQdDFZsyWdfsOmeS8ioxF9MyHhArDYTBNjc2/
dt+kkalBRkPm5VgFGZ0Alt4fy4p6zUm93FgKwziHDwpsIXnjKfGYIDVyWVFAIWsk5BBmN/TqhS8S
p5iYHltTXs7bxxml1/ZFZf+FSGnixd85AiDUsaYD2Ur5KwQylw3GgL7qBLyV7CzRydiYtOpXecdu
M8IdRFMK7bs43MX00FadjkHSLrxbt5LoxDu5uOZzLzmcZwS3a/jKHXwdeMAw3kGlZ1v7TOe7uhxZ
QSa5fhX6jdnAXIBRjmWMVmW71MgYsa5PiAV4gDDw6WabZXCZW8yp2F7QJbLndUZfy1qWgX1/FT+s
B+giRLkVPmIhKniWam/gY4PhFo9//89JPyNroD178RzJ204IaX5U0M/UOpB6lUYV98OITj3BkVRN
NY8yQFReHRpioINQZNf0qXZroebC3ke2M7thinOGa64/TDKkf2n+Gz+evQYnq9oWWCQkV69cWeUq
UaHJrzYCq1aqFWSjR7YZcRcN537htonD+HW7CKbZ/M6ITqP8NJEGnzsmnq5pZ6y2BOfKmL3Lzg4B
MJE+UMnFW+4Nyk7tgWyHXxXMmiRGVq7AnH2zxx29jXrlHhs3toKV+WyFehQ+RN8eWpz7xZSsiEGL
dcedG7yASV1KhdkhcN7YeU3ry3UcwR9rfPAswkisVQgRrY8G9tzP7jZiDAbDDf3EeBHH1s87/F2X
VePKsED2uN+SZrRqEJuQwT8s/1ZjhQcnIZ6QILLLZzTdKRYsLE0VEmPjH3E6ezhQv3x004i2pVka
eHHZvONBhOKovHrimwgEWZNCjSJSBMNtyeFk/dMwVTBsAjAfaZe1psyxSnRiePx6E1dqW/1zSeHV
LrAVoStNGo1Bm6nhGTMey0VrNBBF5fhyGapzQa6RG7ZkSz/jEDIlKYYkoe5eIsqA2eYry4VBy4NI
Sfvxtkh+mQwbstPlUM/DK3WwCXyf2j1LrdbRY0ow2BFjfg+kRNqHGyeM4ePYt8TRyBHYdVOAoE7b
i5S5sxaOJet4P2UqauW4xJt1pERySHHNu3mnx9ngaMUv/vEFVxw0FBvEkAv8yQcDZo6N0ysOHtMQ
/NQ3tl+W7Dt0Z/s3cNsKhdePBt8oagKIjbUkJyPeaPnwXOeF3TUIxHq0B1Lj9wUYgJLfS4mgn4DB
Z8d/xaHSpaGeuynBQoIqxIiLCcyklGlKSrN2S5fjBGb8CbQcFC4b0AO8Ot1xNoQn984AaGWZNT7h
wDBYsmmOqvMagPNJAMhCo61nvvPxKsapU7cWLi1HIRgzoKz6PLAuoTYRHnXCM5SZG2G8CWv1pIp5
xDP8pDPT3e/Ys5thP2WCsv4YftJqu+Q8PB57wTdqxQ3HIdCLwfr3hQPYBpJU9necEB6iUTKNGKM+
EkgM9WsL7e7xRzTG/kTKqZ1f32zuirT6yUaD+xx6v5gMjY56XmxoK1OyBeVEIPALX6niR00GHNQA
Ti1fcNSs/QwOGNTlwnN6E1QsJvo4mTMuw5bMeBMq8eX3nWj+p4GF1vZP7T2B34vq2xgKlDt6oDdQ
SW5R3bseBCt60cgQekcS8kVU+7JtDuv7A7eUCyIMHYPpsVUGZCXf1Gz0dIGOQZRy9SOtSivP+v7b
w8vlyep48fQEQtp+WsPQsGs8f63xffRlcG64StcMy9CrI26XaQLzzHjTGdXReBI73WtsHyvUWnw5
0ghFc9pTbA0tqzlkUfXuz08Q0YY6slr6GevqZzojqH355JWRUAMWu6YHA3fCOpfPL+FAuX6KqcZi
tjwIN/c2/Cn3M0+XZdyaZJtjxcHv9quyUXG5bAv+5jJ3Quw+inruY5V4xqiHa3OiT/9r5uBgvfqa
OOUMyUvEkd6UvCgX+UFs52qhUgt4BmFPd0pE5zzFfr2KYaTuqfxWRAp6FgdeevVVmeU+bvYLCbEr
WuHuwATcAdk0ZqK8Tebjc82euAyd4/s9kImdH2UjKCjtuygL8hVsaUqOsoOhXmeRn81l8FQcMePz
S/Lp80TKAFGaU/OpVhL2vbIfFx5cRBHPxDSpF3mJZy6pp5a7eTphknCvWPsavX82Wk6Ait3Lyapu
8A61bDKJipRP/69acck14Z5JIdNJO2RrmJf9+aaR/qNenh9/9XJoLbuuUcQgFcCPPtJ+pJpkPxUW
dMJnXuo0giLrK0a7I2mOkr8sa609qJAgrNLq79Uz7SSCRAK0+PqpwhcoXdec7Fjrb7okp4KPV5UE
F6LBRkPXrWEW5cgAWIu2IzSn/UwAJl9BLePSX3A+JCSke6a2eF2QI5KeYxUxmbE0SKOMkNVST8al
GbHcXsjycqRkn+zaWvktYEIc3z45NIzwUkh/ffeXr3VGh4ccqQfoNmhlk3knHOy+kyTKK0s39o7x
4IhrxFPFS5AaWNeZqNfzW94O84H7AnlL+ntz8BZ6jrobiNmSeZVrV3/TGI80kwH8phMqyeRKQ9kd
aRwYq5cOcV46sZh7tBgupULpYuozG5nq4LZgwUtuLlqkoxqw3yCoQSTsC8GP3/HX3NJsnPHzSVeh
BtpKxUkHaMEtWsyCayY/TQuAb/qlk+ahG2p0UWYaM9x64fjys72Ee9i8zkdx8SetKxQHxpbmWbyo
YawBJSmgR6UCR25D0aceJMIyasG0l6Bxnr3ZJVDl9/1wGCt8npHhqhY7EJBQp16Kn+NNZOWkmps1
R5kL8zdz9oVG9onH9wHQugRlowia1KBJn1VDUIO7pHQIW6wxWbUq7qMvnutncDTG+IJYX2slO0bH
c9f8ZomiEXzutdE6zBpUU1wVwZrEgtZqwJ8MBTbW/5I7NNz7nO0+WYSsAa6WygMFLbAp8RNwKxzm
UqHWCB//f7cmA0HsAjLXI1au67SZAZxEQ7pdMQb4xHLueeNWP7fhqSpZehXOk8ziEW6QMuI4GJ6B
jEGdRN2GZbiBOFKdRyZWo2YtMYRRWuIUaHhksFluAIvooAjVi+mjOkGCEWVLRMxNfhUjD7InC9n2
EM5NiX/++VZlPS1WFvskOecUWS/vEQMUEgKA/35NMw1kmSlvjd/IaXOFgwYR5D9e2cp4vG6QoZFq
pihAyNTWzkVQcw6dgIntD0x/+4KuBPJClBdMHQ3JjDYHwkdJeRuaX4Rglu5wEyuK35K/o3WwCWQk
PhwyUBndNjzjuDGUZxd5VX9UOpujJ+HTev+ictyWhKB1GSyL2tvODUWW+MvwWn5rchw0p23EryZW
WdnN8Cwn615QtTGjBT3xdYM/S70H+ITbwpo8kOkaJkVOdozx7gx3XayTnsRy+6V2UgpJVmH0rqD5
wTfBjX74yuA4CUyA7c6wKQuXag03mXMWaYwM1KAulQivkHWr6wyCOlHRNbUxJ4ekjNe+uxkusKOn
YhrStkCb0GT59RKzA39dj9lO4QqdYSDrrNMu/wkTQc6IQ1uJBdgxlk8Zmt1uCsTRxrtwQk1b9iYq
bqItlTIqZ02y9GsQegIr4/+/vFelRV92AE+cet4hzRXj8tOMS30YIVFnzfQD2qhYopw75O4HagFj
ew/L9PGXhd+Kcwuk3bUqQOKeJse3DTIQAHRl8C8Y1GNnzPF7ad0DUoaNdf4w6oc4IbkXM8cmtEcl
Zs/1Ih4di00DoR7jy62tN50Toj0ByKTllyJFsCEZrGUA52Ta/by4FcrrQrwT/AY5DXMQuHelARY9
6pgALVatyFezRBlfm/yl12koMeKM2PinzA0BWQOkcEVjwMFzKQ47WWSwiSkdq1gC9x4ZYkcWVE10
bcESNhu4AwsDcMzvKKDVWFR0tY6YDOc+kuikJCHaRFl5mHNJc1mJC9iZScG3jV+2i60pG3TZv2rX
wZEqJJd2Xs+V5hOYdzNfIf7WNCC4SffnVUS6vwvKaSTn6sCkeXWDQtcsRYEUVcqph/sK2m3nIwjz
PU/bajc2xaHZ9PhUm049dFmwjHZpXseU93fu8CXsTEf32q1Kxs3pshasFP4r28dsOmZsaco8jqe1
PPOEKKc6Pxb1veGV9qIpkl38zHOsBwgOzh5BRMaW3nd2f9AGKNmLfeZA5oEhsoP6m6/pCXZQHMNg
Vb1OfmTZrhsxAJgi1P6RqEvKGvOrSnDV8By58+qwY93xPQw7BnFvTqZQ8EkpPcfBFz3Vf4Egqb5V
mzRhAwyGI4Tf7IFfyaSCxy0ZtAHNrELoU287ljByE7+Elmd7nNGuOJGWjlmhCoZLbm16c6zS+yCr
JRX8ygf2VSQtulAD/vyg93wDYZ+uoSsDJ4iR6lOK7fKRmuOa80xexT4B1KIHVyqcHD4dZExfG7WQ
ru2CEDlAxxTTiw2tFUkPd9hvI/GwgPRFxEk0teyNk5+XsmxGr/+jVVxgBJlwj0eKxh9xXfuxA/a/
2LokQc9onhiausl9CsbzVxqzZJCZpr7JOMVoLQLNTMqEw4NUVVg0QJ3580qiIhynCfQtbCC6+tFI
03T6HkJewruF3VZRl2VhlOR0dlfAaF6VoTzg3bBNKr3VOZ9Apx84lW3AsVzFkFhHinc5j/ViV353
tGJlvE/JXB3uC5WfcathVupvo1P10BVWoPzmoGtu0B+L4qRF8AbeXFQy5rHYK/m7XLKjLj/C8+mO
dTQ4t4PnfYFoeeqcZgunB/3hw4k5k11k/6vZ2R1ziIS4YK4atnWtXWarnSsCatsbXvE/JtwCQAAd
A6dUZUKtUjU8JxYyTCloWdSxq1x+4oYFA7lQURelFuV2KmVKUQAz2MNanz2d/J05C8T3vR7/fRPY
KZoJcXjxIEbVimKSBQapOKVurIW0ug1G2bLlQDuYopkGbDcGfAWY+at2obllo5DZ7EcUUSRKTooe
LC+mywgJLuwWr8c0eDop7Vn8wIZ/+Ve4UHcpWqFbbZaEkSNQ1iMI1tgG1CK14k1Wm5/gxyqJtRCM
rLA2T0hYT4ml5TteACr8ISXeZMEFvpu5QBSlIrHws/9PlNMQlMQ3c50NsEw5kDK2gvuhpb96YOMf
05LvLrtbIFeeEe47iYHFUry6MSbyrV33PKf5bLboOfhh/q+l3biukzvBfi6nU4h5d9iJnMrluRSY
aP/7QzbHL0zi4KyNknz5vCaj91WOnIY2lgwHn+/EWIK9du4fs1TX9WIGoUa9idzJLkw6dqY7i1EY
vA4QO9avxcxKsRlF6NSqfQjSktt3R4baI/MvSeHBVrYjgmLokEz+4DoSnQ1RSkhFuECrj9nBfGhK
fZP8eE5gaCXQ+O20YpzcNV139RkM+xlk6Iwyofsgxqo2WUt3InjxrOoJZNtOc+qqVEVyA9SHnZEY
Aia0TXwVAv7GJHnJnMJpms/VM7S4+o2Q4wZkC/nHYPAZGKsLavN6drrJyeYCVAAx73CSaY/EyJu+
jjrxQvgV1i0DTtwugF3l6ZKtwmlo1QrQIVj6i/f8v/RCtmUUPFm7f/ROI+efxNCc8QF8zm1ymAJG
OvcYBx/b09/49Lp3xskB6c3SdVR+41VG4KkOJT88eA769Kqyu5aJQugbVaYI9/cR5mFF4q5TwrE4
qdv7F0+GG8s/4a3b/+F9chZK+IFFvsSqByAbtWbR9B8JknQKSuHC8hnebG3FNFOHfz+spk/OUJ+L
2Elq9IH0t+SEPu0hjWLhV/E8emnH0I3THYHp3p/gamkx3KS4q4mVG5OR0mgPvq3Bk+UWETgJbkWa
YDfGNFJPX3QbSIeft0/h/ee1q/3f3aurzeDWIZQEDoEX6PeFMbprFz2U/7BbdM0Z2foqI/AOsttX
ABO17TB2nujv1TVmCbQ/94vW7/IWsrJ303hR4EDm/RdgBH1wA+Ic/R7MyoeoQN7x7ceGG3FpHSH+
BTI/Ul5rxZIjNE+xChXXIAPHK6t1p/cXxsfFdok0K3CdbJJ7CetzpPwHl1V2xbLItlTf4SyQ40LA
RsfUcpht9/di+RyduUkfaikbHJvmW/A3eseDJWT1TxBp4oMgABuSUPgQm0i25vKDt3vLVdHvYo36
YQIH9JwAVkK4mavmJQCTn9wRFHnwOtjn8rU2bnr05xFRgyvS5ttPLrPV0Pa+oiwaW83cpjONL0NG
8IX89P+PubXctfRL9gs4sp7W2S3TH7Ji14rfOZl74THEabcvxhLeCIXrlwsEh0AY/gHyyRCNA1HZ
sZMfd43YmpiEVIyT4SfyBJ1DU1V//ehIpQhpQSCQkzQH5rbkRTCpvmsQ3tbM09Qt7yL0G6/pY7tC
LGTb3FhMDE93mY4H2P6VJsZotYty474kgHQDK6+B8yFZVGpnFUDMzTm0MZOpi/gl7GsClmbo/c86
gPC+ZAkSkcGdlW3r6vesGOeCZ8jmqmiefVQKJIcr/ObaFQ+n6ydNKKAG1/XzYeANgEu0OviPIwxW
HtClnuYiG0aP2aNcKrbgeqBP32F8wv68LptChXXPV35uF2gS52UpidokJ2dUTS9fuFfJpitrvejf
dtD6gS5Tt9HafqQ84h82j9E/A4+6IoRc46ym/akYjLBNFSSwEqlWjJHELs1dnzLt5nQKyIZuQSZR
MEjPtyZiA9TP2Wueg9NH/Ef2Drak1jKHxg2ddN3nFLRE6QEaDHic8UW4r17RDH4jAJ8G4ZEJqZQu
D9NkpSzm4hPgV5UJjdMFkb+YaXCSUJX7FFU/ssghcdu34Pa0X3i/0ZMLpBQ5plOgjUlrW6/1sWrH
Bdyq3PGjpHOz2A3Qkbhvgj/Xa9/qg0+qVZKTifr6+/pp1saozpQTyWsFpk04t6TkELxeNFmANP4M
H819pqtXOcxS7pnsAX6ZhbWLpFUxrbGLxvAjZl0PcKlUm1RX4qOlAzOqc8ECkPh8wWYb3KWqs71O
oPA9tw//tLpHNJUaagFOwpQ7y0gv/N2QGnVox1ySX4o9R7RM39yWd/ohRyNjSAllnAPrCe7HxT1j
u7bdyWxvFxDxtX3lBLQ8Ks52BbbCyhCWx49LT/luw598kYGwIH2FBwgeSro2H5is4hRGGlpIQ3Gs
FZIWwjjXUuVZv173bSdKDowyWctjRVpdhJ6FSjqHYgdr/YgLZuY3/f49RnNkdHt9a9ipzT+Q/SUR
BxFYAYwtpt2F96cRQL1es8wNv8RV6IQQgmT3ir69iP/jDxFyZ0p+YNHxw2ypiNthS95zePQmjKKK
h0nzYEQ/mA4DQ0oLsl2IRJCJ98ik8T9YHDdMOV7BdBQ089YLIW7+9+V4CsR1npOL+kaDSefVkpwp
nhL7Tw9vUp7I8Rk/GCiqQdK260Y99C5E1mqop/IjRJZIHJ6hhpSSdPgHfYWBajU2Ehda0CP5DOnb
At8YBCIPoHAFdLZiNtVGaNcE+bcCRW1+sJT7TZXXQIp/rElkukIlcsqyKZjVMP1eIeQdj7i0hVYC
ctHupBRrNdwKBBBHHFV38g9nm1lMKiGs6J467Tdg/TLMWwR7MgHJ10zoI0Wd4fmyaK8QyZhhjtTi
3NRfccPr1cgvjL56QNpCZfpi0/gRphcuz8eThCiqGVlaaHOmIswfftOfVCsqL/NbSyUdkT7zDqXX
OjTQIgeava6l0/ppR9TfjRDfJWI51T03SdXKugZk/clWKy2MZ7q7qadTJ0xWWNqC2tnXpL+pjrrh
FT+nq/L84LC4J6WKAGYoo8Lrw9IClZ0FgMvxHiageIDqZVjokentFm4GztXzjt3rYg88Wp761Ijk
78EFzeKQ/D7MXOK/ULVLYbPiEVS1iiqyZUox2XrzFGSrrngJLA9K8t+gnHeF9KwLWMvGUANseIPr
pDENI0wFW4lHi2LBjJNx+lIenceSTcVhJfj0xjggSNwsBrNUgHhrqFH16dCe8Dfe9xVU9mT2cG6P
iVsHN7IMajw/5axU+9BAINDFyTpXXNO3HOvgY/Zwg/pjuFIK8siT8IFHpH+O8YrnKCJtiOKZPFoY
Ehu0xyRMDbEL7OdRgAsU+2r05GmJgiKg1iM85SP/FIgL+WnLhe5gnNeWJaWI+JN+iFwI8jY7JXz1
9NLR64enMPfscB7WfQsxwPTP5Tvjl/qNNhDS/aQfCjuKACYed1PGn1sbXtcqp99Sqv9Pqs2EiCX7
9mHAR0tbkBl1xb9vJ7QdGu03xRFoceM1pEwqhKfQyw5TQfadgSZaAnmdtlUhF1oPFN72l9P1sW7p
3hhcayggHf74HOq402BulY5kpD6PacNU73OKZBXnjszm0TdjnUBU74Ia9WeIQBU4SmoQho6gWpbR
r0hheo/EZb27zRh9hXOjg7d0sQBaFPitDzD7xIu90uLqFSUTmThTKhKqCaZE3ZXcPPSTvkACJn8c
KdDIcK9vzezagt7OmGe6Ed1piA3k9aLCLOuaj3YoObWudxaK2wA2zI43+G7haRTjLv0t/z/E6AxW
krMoFToREwWsHWSHfVC3aKQwZIV3MirO0+ua6VWJNDLYYJEKYrpujRGWElcSybPs2WRxVCqK6Hdd
6d8lrEWfZQzshetjEOytZpvgRq+VF6pjpMyVHQHw8XZl4QfMG3QmqT2/NVHydTAS/JDReDrUY2Ln
PIAbY8cZr4+HIsuHZqPGN+ZXRI3tDZHOlbi771BlkgaEq1CXNGin0iVGwxcJGI3KxgyelkmbZLYe
WDdQNTRhjlDzIm9qVT6KXez1bK4YLHGeEe2Ev2Gt4V4HZEjpj0EUrubGyOMLWlMk/VaOiF0zlfIY
h9zfagKS2IYnHwpGzQj4UQ1TfD6odipSawwB+BZvqQfawRiZVvTKq9XVg76v2GpT63RO2g0qE1An
VEcovCV6NUGV5eLXAVkVuVgB4s46o/DnIsUnu83yI3wuQcPsDUYPCCKYY13VBcLF2bqf2NUJMQh9
JbMmWn/w5QHH/iseh4wRXZD3fS494AB70fLu1kP/duXUi5eMsm6n29PwYXIYBteMLS7epMfplSq6
PqwbVRQ7KNl4c9EJaqW5ZoYrdmrqpb8QzXwK5Fqtm5EsSHf6TajDtd8FeiQQU1w5soa5iZtozqxB
3Gy5/odui4PfHKhmTe0SHwgVaWffmnpFoVdJxZbpjVdP6Rg7YfkaPnU+y6QJ0HVP+vXVdthbHxIZ
Gk91iKZ4G6SW5ifJ/DpRXADXKDwY9OejMrVTUQGhfaU0/MabUlErvnXiCWnlKjWwiPuTT4ygYXRX
n/Lmt+WmAi/ZOKBX03u2+UXzNHif46tMV3esUTHSBLYuA2tpRNGHYOkbHiEqMyenaBxGxTE3HUu9
QCfyiwKO5wcRUHj9TVhhB3BaqDe+ikc6+Co36v3V9oZl7HUrk8rTi9PA23WiHO2vXfjcVBsdOavw
S1s3iXo8b8k+X4JhfpZAQRafeImZM8iaZldmQ9V3Vy5p0H7mln2NZTx51SkwmkZw5qh9YJx0DhZk
/D6C4e5Ry8AlCHuSMp3b7ytcCTVUM7SCEOgoNKds5BzkoLzqqCdtXv/GYhE1D7TBnNtM3/rTpmsl
5zh5ZYCXcvNDRMiTDo8d558jiq/EmQkdWn+h7Rg7sKYL2sFqKKj2Wcv9IwhMl6cFwjJKfLJHqNfX
x7/rScakr7apUUyr9R81GPLzOlNQqPH2NUjDMi4IBIqK+GXYP5Ca4fk1maAVMXk1v/VX3a+BSZrl
A0dav2smAqy1mdQIRfDsao6KxP/L6pN+E9Ne1SOAtEyS3X9zT/uEvSIs+ECD2FcywDfZS5UzLY6/
zDTaSNUF/i/r2h8km+heoM3PwyJO9TV4FQQaSunUTrcCm1OjXummcx9wZAqnF/j7R79Cq9QUnqLQ
zSK5XhuSrrsRDpXjphcRKZY1db0vdc0BX3Gq4O+24/sIQr9S46JuWlpOaAq3GI4kMU7Bn4O7hZxV
k43AB6LNJ4fSBNB6Y5TOU7jNKYmaYUYDlSqQts1eoj9SjGp6tJoquLcz5SXyBU8i9lMcyaqT1tJU
BSdXYcNM4AgyAVT/U3jRsuqLa2VbFHvMcgyTC0jrYV8Yj0Kdna9rNMJ0WiMUFtaNGqCgvUC/hqIg
ij7CrfdmuZTmUIGm+FvN4JscmS0vtr3z4vKa11H6PrWCsYlQDWDVBaiT+fy2Z0NuTteWZJcXPYjO
thy53LKcYucrHiFNApuneil5hiE0hAqVJvKv3N7jCmTDsBQM9y3XPQiI3axSIAQb0TDZgTLNy+Br
Qm2dvoC24CMRFA2YjPVgGsGJaGcRqYN9VlA+iBQ7H4x9rF/pouH40lfYDjuYbSZyuDutqrG2QbVx
d0cz+H5RQfie0kUyfBanpFYgtk2nBE/NTPlmr3Zwit52RI++noQP7sEN1jM0mmae4qbBbvReGgA/
H9x2/LfG4fEOmBHTTGsAAtLhTmIZ8HGzDz8Ig+gKyF0kh9D9gccTG1kesjETrQinTfXT3G+/zL1+
At4ZlaXurMjLN3Cn8kP0DT7ufI/2LuzMVIXcsk55fAs7YwSoQ5tvpQLIB1Gv+HC1vQHLTmvJ1stb
Wg1msI2e7iCa9rkstabhUbRjUkAB4vXQo5t/8ksGrdbn1zm8zB8FV2uM01axnXoQAFoy1qzT0dTo
VmeeHiQD75otpgE39fjs5sTvoz9L+yOaFVmHCp7IYT8XSB6/Yb0SIlsXbfbND5BM+FcQGjJRnABa
kSbVTR9odcAujyUSqdGxsdwWaOTqk3VFzeSLoHJSUHCsz9Wz5y3NPb8SOwOXOedVAZ/4GDaRvi97
TeKLnTrQdMO5HhaXC2WhKzgfwvlU68+G7HdS2lUI7L8UchKGpGe6rb8zQ6UYYTcmvK+KTw0k0b83
DzBoAMrLRVVro8pV/JpZ/YdvYHyIMlRdny10hEGzTYJFF6DwTBw+3aREiGu1z5Fj+NPPPUSurdnN
a8c5w8JTpcjHtlNMn2/I4yximb5ZWy9+HI0Ipp1vsmuC/wHcfLfRJdaye84TX3mKXG919ThzIRQT
lKHZzURkuhnVaOpEWiGEWKPJNJY2ixreWS31yK4N110E4/dHNsdqzazReKBv+nD6sglIKbgUj422
0jAiNJFkF1QRJEE3L4TpR3G3VPs1aTe5rJF8fkKHEUTfvm81QU4Td2F3hbg9fTuhWupBZUEdShRM
EMUm1oqnKbu62M0sdOIdigcbj8LOJHcZdnyFkFXMG6gFMx+aZQUcdjg2LGONbrtTUQVLGkF5aiBx
u8sTMo8NGaQeED/z/n3hBfKtU2K6xzvYYb/f3GS/cUzhJzEXSFpAJx+O8bGnX3Xv7ke7BAU5WLYx
ok1NQ42D2C6JJu9VqS/o/M3RyHBGRTHCC/IVTtlk3XLYgjyzLcnOnaLqPEaf4vba4r7THYeWEuWP
K3WktVvguuKDkT1uww2oHcPLFToqSCFRiFOvDh/IeOHzw/69PWLqXAR3fYvPImfZGdWk76lZ18FX
lS25s4QeUSoZvmhkxJOp+voNBTVoCcJ/k40gcKsVYjPChO3Y9KBHIfljwQDfy2e37DublGBHsOC9
AQPDo1KimqIGGoK05ZGvmiG/D8w7PU0AWoZ7m2l4avJhwiIzHoicUtAugwwk0DXGPuvhhpNGLubf
53mvr1sBGQFK2bdAK5mh7ZaQW7oOM3mqlsQtUYeMVpnwgdcVYRvxqC6senVPKwkcyFK53RXKr87r
Yux93OUe2ns7TEcylUpplhNNhmDDitrvZHM0vwsT/IaJA/LS2qIZenZ0iHV7yVYBqaTWudjbrQxu
LrIY8jozK6ZQSTYgQFlFklL2xTTjRGQndz6dAujIZ3O+aTvRyAcnJ3TB+icf+a6g9cftB3/6exgT
RUBzFH13mpYq1Mzd49Lp1un7G4NNJsaibXH25yKbgUMDoh7onh1C85VpYxbUNnROrDpckjASRWNw
aAPBtuMNlRVqrdlFijCI+roGHJbnk1p/bSVEaPms1vPMrOigMjg7gJH764BrRZFtlXJN/1rsVLoV
B2UuUEOzkpF1fD+gYbX+MsvwWMzOmufTzhxf+/4e48KcyXCx2RTjjccif7CeyHt0eBbtJ0wJAJn5
i2XK2VZ71302fTvlRuPJTurfj/GmqibofgQ+xjzoeYg4KgFKsQ3wO1zweBC5ZKMN2TrwPaOQ4Mh/
1IUKtxHjO71yMu89rdjU9l8pr58t+K0qCTDjeg8ssCmPUN1iV2H7gpJ3OHmFUQs9wTm6FDzRWY5p
pVfN3xV9M+ffiLyZc0ZYC2TTszpDHiCMF5pO6YHwF3Vj2bCYWrCprgG8A2+1vVAFS5HFKMKSNYmt
c7lJilnlilBabDtpoKvSZxlcN1GwISHv4lSRhlj2zR+v2ORLkEvJ7/l1plcrl8O40UakVMTVmQL3
XtiBAO5qoWz489a9j6zbv7P72AbLHg7sL0GqPgUxmMufOIDvgRJN+9v7hsjJS8Ai0+RFps4P9o5A
fjiJYyZLD7AZgYApRENav09EL34JnPbKYP2wZggNoPNNLELonpA125itht5/8/4Pr8uIPnqPBYWs
bRn8eo2UMvns/RRb+gK3i3OfIVV2XQnB07Rnf4v89YN2S/+nQHPZSgTaLjkwlitGjdQvmIOY7hfq
ECrQuNNAuJ8Rlg58XFwZsjIPftR5vVyBRDx6gKfqqQs2YvTvJhp3afZRYV9yxEd7TTXYTFKeYE6B
F2nVPJX9MDKHf/KDmeVAQ+yeyPVki4UPQs/s9hT4szyNE0SElviSazAkWhYtItRVGhJ3h3sw0hIG
p8fV+x3qdLmelTYECWoMw1Ve0ld8K6iQEHuBqbsPO/qGQu3BVjFHsqy1rU1/gpcUdsGLXV+i/8d4
SBnOSxWLVRtknwgxt/ESwuIVQ4yzskqAGdS1pzuom0LMwDXRiYJQCZO8Ya5vYbTiL3vmns1dai+J
a/CRwDDdbYz0M+wmO1zaZMV3M6pNzQAz6o4bkM/4Pk8kuwPNan+Ri906y+1S0crRyQ6LyS3+rpQX
yiQKNzT96TJmzX/SGO+CfBDYQi1yO4GDAyiSjQJGYIX7rih1qlqFMrTyCxD/yR0F8GCc7x47QXIT
s5aCt0zshB3lYL8Rv0/XwGdloQ7ApBk/ZGsM5K3UaKVJ7Uf+jjn6qQKXQMSq4uOuC1waUSUhjqdQ
AbnGycVVRVAc0EK3yJC/Zgjcx2EAZD+ED3bhH8pn/UON8gFr6dN6M5wuehruW7RD8lhs3xWy2Cju
/I6mTN/YTkDhTflqDbNv2vLXS6ncSgnjQezblxQrnywpWlhKTyMXO8ZNTX/4VZvv+7CSJsnPp80M
LaTyWnZwhPCSSNbKaLjF1HPPyF9OtmVhQPUzsV09n2jRp0SJSFapb4ctY4Ug9uA7Oni3oe0oCfTH
Ifl2R4fGPG/M8ZpmUGuxGTyvy9qim3p5aJH8RTKsD9cBTQhyuLhtoY6JRRhZZq2xetkKj4SPZrOJ
7gvawOQmvrwinPTEB/gYJIZ2wvZ/uURL0WLb/FiLMA/NelXumWq7+tZHkP1ZquRnuU6qRGs+Qg/x
8j8l1thhJp6Sm9FzwRuRKK3xtJISZXt2uwGBkDjnMZWK7WlgTOI1Kaz0oZ6iyD1gutTSy2qjzAuU
Ih1FLllvFYBiKYf4GKQ5xdy2KsJeZ4Vw0zbz7oqv8G4G8MRxAPEhbNkpAOyYRltccIaTDbxf5o2S
q29G3ucHwxG+Mtc0YBKxcNU1euk2ZZXO3Mrz0W4Nw6QctLPB5Ud84zd4Gw2tfm0FXB8O8MF9GQ51
V6w2hR00+8Qh13rTPDskA8FdnOqyVkRc/1GOBv2vFH+ur3Do+V4QOU1LJPOm4FxJuRTJzHGe/9D4
+4bi9oPV5PKFEVtCnRu0Ephz7LV0QnOG+MN7wCOnzHiO+oR+Rhrex04Hy9lA6ZVWUyignArzwhXb
nBX0oAcK0jnyxiETvm75YFLsvCrGliOG9Av3OKil9SuNswFj1iIuyxW3/KTkqt187dCDiVPmrFn0
YPryyls6WV3Lpw084kgli0BI9rDvlqKiQ2JaufFXnQoAWgS3zSgxQdSSXER0lzBFweIFNkh313EZ
v0Fx9Ad8Jg7qeQT/wOtmzMPwI2A9PSFLVDKyR802Z8wmIN662y/fpaZlHF5HNybZuWuXFbJhVNvH
TGsvK1zuos2AnXSPG1q6J7NH2VT4lk/5XKDPP5W6iVHCdcZCbiyTvkFAeAymhemuZoiEoh2dbEei
HPBzVDTaHxB6tsVZTrfg9tWxXNgdMB25/zsG14vndWUUYBHszI2betinIQEZaFE+BMXeRkkmTl+5
9AJ995dEIETKcvXEb6JIgzMz7f1NZLNPCbYmJFgW4K25bs6KQqrIZfwvnPmuoqnKUlE8yYu2qv2l
UBwTLWERewcnSBOPRwy8iMimTXJyLl65mSdtYUJs+GO7WG8zhu4x6BQfpgjCbSOISY4XR5xyLhXY
LEqcte31/F30Tfld9MbB0sfVL5NuiSkcB7XYabo9tV8q4JkmY3PgkTG4MqIYDaqEwYfHLj6K+AkE
W9kRaw8IpAYSyD2uvmt45jqtAwVCgShXr52uRbUBgA+Z/68gFOtRg/7ucHIr9A2fO2s6TpVMSIFm
5i0YLeWsqknpbCmzhfS/9mtuGc6RWy8R77MuQDJY+zcaNDEBma5zf0FUMF2LZWFwOz9Y2p/b3llR
LWUQriN2sjJ48RLO8V2o+b+BbZrgykJZyQJt7/L4/dPZTv3j96K8c1biq2WUEWJ7u+B/VC1FcKX7
nXRZsXWluLYodFzdtCe2mDF2JdHPYgQh955MkhYYeVa66mY8vwtwTCIAdFLOHnAYG31UnoVWIXtb
pB7pG90Gl9xyA2OtjRlgQwGqWaCxbLsvTO3NN9omOk/hL+lme1euYdLqDb7pVv17mjXeGIYa+eUi
8/l+VEdc8RP0q909cGje8l6caqQ9IvNLq8Jg9Cv8arE8umilfo2JLrOD06QfIS1mCuyWgE7KuTIn
osDJlbEjurgQyzEC1hkD5as6gR0jCIl7GXz8X7uBW858fq33VM4AFJi4BQiGyyWjsVrL68yOYtZk
zZluoItD1JhrFl5tDrWcx+gNLPtxqB3R+lLBoml/tWQeQKUbvKchqcdl8iLUsoLlrvAO83aywi82
pspT3lBj76yHZdGLaqeyuwtSbCudxBtusmTF/bNwXKRIxcwKCjl1WiS5AX4crJC+CiSw8khsDYOF
Jpe8ohKCPIeGd0rPEdLzCak9GpILyN5zHUyQJxFNJqNft/P/ptI2DYZ+XS4k4OcObpsetsJOSJVZ
LxTQUD2OZACR56iL+tjKdppfilS8YdH83uqXfTvzoiW7vFOZGBi5LJYLJWgiu5DlMuM/sXu4Cdae
BZGWUFvwVLPcgNNJTwRgwL3xccBAWaO/BKT4pzlsd0SE4ujlb8S2E41gh/9U/YED9tCvoSzzdAAV
r3ZgWrio357tp6Od23/x3538/t2j0BSfIC5KifVY1KGbCrYAbiZ6rCRAWumOWCoJc2H7Drh8kb0C
1DTFSvQg4ppDUHzSVetYDgPDpLtlUsd7/xwNkXx7rR9kyMwpVeyPoaIGJQnLzFld3m6axLhVncah
ZSMzWWSMHKSNP5IH85mfGha5ahdaunQ79CUoYpLChteWy9rxaG6tHPGmAMS8wDHjmxafYVv27eHK
8QLk07TxCg3UvXIuHoePpO1lhs09wfez9SRtAsJNIfzWeLBYNLy6pQhtazhUqTeYpGI+tL87QpSn
9o52f0A/rQMSkydXEKiK9ogWYIQukIqoy/jISsgtrAZiFTkUWgNoqq7t64nFqkuz5Ea5FGXgsHuW
MTL0cAVZ7Ejz424x9wJ1t4e/3a8CgzG5HQfhpJygoWzta+zFHxc5JGEilDauz+jq/J8jLoEkCngx
zZtecUy/pftsq9JtbCWgFjgfcp9M2P3mDGKpK1hPxx9F5m0wjFK80h432jYM4qf2nUHlb53C2ofH
gwbtVs3ScX2VhEugu/tGxvrf7Ac0MXwkhcddp8N6WxMEd/8m/qclkuZ+/7kl75shrOBJPd+jEeqr
2n3m1d/jqEFOz8R5hRh0HNu29VCLZMf/c2/9kAg0FQqKWttwGupSuAmutZNwbaHi3UKJvQ/p0kNG
Qm0C0eE3s/3z9ZffB9q2JH9Txnfv6cUgkeMUe1itzNExuM3aaNz9t1Hg1NKjsyCihlLv5a8aMKGK
fPaygYq2WF7TzdcsVJTOp3/zc2IzZcdsYJyuYYys6TOAEvBRcqbqqAvkdk1lMATvklRE7/cancji
Fjb88NSHBgL5CqBRqEN8DoTYIu/zwv7aXQ5z7mzWMq1UnjTfNVP4fmzusZA7HYV0a2AFQZk/rel9
oGWXPGt+1ITgBM4wSUgYZ6RmwiSq3jXXgRGsalEUnSxHFLfVD2Q0s19vY7ze3OzhNjiQxDMOnovn
tEMtbjyTDipZVbw72trWxQQcQl5XAGGJacuuw30aSP8AWUj0rCK5z78O/p16lgLhLDrubZ/0cwKe
xWngnO/yrOs1FK/7cEJElLUifkDG0tQGobE6d/NuciFtzLmCss6Lc/0RdOKTRRstleFzJd5BjGmp
KNCUQiF//V+p8M9kMc4x6Ldv9izuYpn8bDQClZjmclLy69c+rQ7bVyDyATYwazwgBNN6PM3fm++o
1Hm5hLmO8coWMjVud41x/hviqkJrWLbTv3XUrQWtuRa8yGcNa0akWdnYiQ0JaI2kHEFHRONAXLvD
PWfW3kMMZCgHbfb3SNgyMT/u/1uTUnuALO9dAsWG0mSvadI5iK3qz6Hs8jpGpql9NM2SSG2KNnaw
7+QmuJEkIqxCPlutIIebyxRiEosZL7dJfb6OmS4UqytAW/FbcNTbH6BYZdyMA1I322l0ErwZClwl
Q6jQoKyezXoKp5vvxTMHk6aZGQ+xYUM9E6a636i6fBzkHf6ypR6oSLq8Y5er0I7EdDD1PjLJjb0t
stsUUDKDA+uBlIzF79NVBHLcAOd5KHF+U5VMPLaP2PCGMRR/AhoEwpTHSUoyojUTo/tljchuyNqx
DKrnWdWyUHNZFac04guWF4csfa5sYJhNrXKwTQQq+fci3/Alm7pV3mfgN2TXLEFXuOHXQqINmGxn
i6/wNJLG3qAOW6rhntzzsfVnMhvDQZvo7iubcQ20E5V4FTuvqpVT8tnqCsVtyuoPp5tZdfHnsIxG
PLPAciZG+xsvjwk/PVbohJDnuf3kV/D64dthDlQcczQnn56thyZQVBYAvRHpiXHtirKvo6ovdz7p
XXM9j/ZJ8h6a310xCNud4rdrrv4M0zIhvmKBd4tzaTHKhnwGi1JIMuDoSYkp55mBdyzsIuX/WztQ
0YluhIAguhkH0nxzlmFaDNSbUXf1iZLV10wVz+Ma8qBlv5nkDCjOGovIMO4vf+/F45uJxSOtMPOX
tO4Q2WuWHto8TJLFcvJRKE5aajkgG/J6F4UvOHXNMT68PCoNRHYz+IjyEVSVQBWx0evKeup378ZU
W3w0JlDpPkVlqn39VbufFo1CK62t1yLq9RMbwtc0dZscaUvQHVjdqqPe2f075Mo/VP7dKEfTm9Sn
alTsopl38EVHlXDigK7dXCa0HyHbyZM2vOT6U4gtpz9LK+9MvD29QnFtpUKrEygDWoz7vX7RdBFQ
8aU5TDYE3Zfseon09CMb9cAHnrlR8M5hBQ8fqndwSoZms71F6oJ0gd+WSsxXhxql7JB1McPvUH2y
ljPVz1NA660qmM1UrLLYjdaYJHbpht9hjyEOp2+Iv0BQT8oQpqiOp5OszaWD3vyhJp6PXmzN7zsa
GAR7/X1uIWGN5wmM3x0dR5Utx0y7LTXZrHEWalAlx9s3WGFPiwLkXxa5XMaLOCyxAfcXcHWP6f7V
HvSY8MBKXhgR61IPPCUePKB2Ag5jNFOCdV0tgFt7OmEpJs/eVXdFF4kw5pCLRtw2xBBHEWCdU0Aq
UKX9QLqtpiro9PKi8vRv9K+UAVLd2ygw28SW62uOgL9mykNr73bE0jtE1IKeIAr6mX33wdF6VYQs
a/VRFNvMhCXztYZoIT67xM+YxnCtMTk7lpJWFCAGttot4Fth8ntOQlbgh/mYJQbApz2y5eWNWfTi
5rA9OkDCuqI8KK6x9gjPdJtwwBDV/F+Yh3QalhiCwQKdUzJimewp3iSMrClsCelqCPZ/eMhDHOLd
sIEV4VLuuHfHlwBF8YNGUZMpElNcI7cYLhhsn4awMEF4tJ4yq4hTenDQ6G2oY162HjQRceQIzjgg
pxGX3SiDeWwSA7vsPgKMCGyY5Uxk3RaCXes5rR52hoMvtl4pS92W75MgeMqzg99zP0wx96jUJgDD
BDCY/ixxIvAETgQ1DetE/3EOAzNz2Zj3/Qr536ZIgHrmWtc/jGt4irDvsCQ4NSpEtgs/5ZiOqhoh
WYn3SANnWXsGk4ZLaPQNhJPmsaAX8FBp+8zV+musT+7jbivW5pGKxsFK4O5Xi7pUGmgHrlI4uwFi
ALOWr1KTZGf1we4cYPf7++Lg9HsOgX50ypvgqE1RTIaQmdjvwjJjaQNwZcOncWzlvHWRo28SYdxs
6dRCmTFvI9umAjOTDF39dAjBwKb0S9xygJ9dcKmyUYXYUW8tkEykw/+huv0AMhddVPde/L2kO9Hl
1EtteoU2Oug2QuIr6m73ARPsQ83HydNOZMRtCHkSdPfIdI0cYKEyi69y8kLBdpUFVIXVelA2Unsw
S6NQnFf2uxhCVqJCno0vVhxNhWrhs9Vstd6Bvhj1V/JIg2OsmL2o7xg+HmLY1IQJJb2TC37dvV/K
CoIlM6rE5tk9oYKexBjYok0NXtA6jrExCUIRSZEQ+VUlt9qu6GjXM8JfoWkONwRJanjl2tMiPi90
wzihPzBj952U4nqaEDEG31XylPh6w2ke3JmWiwn4VUD2RRWsiCeFQ7tX0TpFx8meS9ssbTfv7v+C
tNjOljbCnU98+Yip5NFlI4KFFNfZxIF8pwz0BlcXvgL1DxmB6MOJTMaelvfnYycjZUeFGKL70wdF
/cGrNc+GJBVe80s+or/mSKwnVS15ytjV7WTSe8uIPzDdV6/bRcCabAaQ0dGebZSB+WvBnWGA0TGx
SfkKtktx8BvZbUipi/Okq9Gch40yOi7sguMWhwxWMtc3ssjbCHvi0iYJSEXD/2NTDNNQGCP6V7T0
y6Jxglco2oXQoF5w4gk1LH22nQxNOYG84r7qrIANVpLVcIxB1O+ydUFOa3ENAi6PlK8oDdP4WtVR
KW3Crd8FpZjKzWv653f6F/naojFZ7hfTWdGv+kUSoT/qTF4E5C3upUvobsDh4qu/Jv/mvEQzrH3S
eRvXx3Inrmh9oi4ndRyh2HvrqPJbk3FxGX7y6BR16o10AoZM2JKLqi2chOWAhREtQpn+ytamzM4S
Rtc/a1qlBHkcmUiAox8jN4c7yPd0hmVhV3BJHkqOfBaAYTOdebgXdF02WWC1yHdtPp32zTtDCoFl
e7H7bIG0D/vCMEj2yRsCBFFB9l1+Q2tPknHw18EMptdE8u+97XEBCHf/DuxlEpNfryW+q5tq3C0f
ja0k1v0M80dXzK1eOzcNTMm+sZChfXbYQbebrQTHXdj9GolkKM6Rx3pjBQmWFzXbnNfyDZ04mjjk
yhc0kFmpU3JMwtEhjbnLeJO3sOcuM5+Oxdjk7vS/dIe4tWSIuecIy32RTmC4ZE0moM/uzGW9SPS4
R/KKQS99Wzp+rn4lvjvpUsGNr82l5g1agqYoZrUw+rh83koVi+0fnuA1odPYadArBABgj0TQ7Quc
/aLMMYQMb/5O9gfzl4x9SmkoK7886XUu43aBALKvJw9+IKIUwvdqwPEwPRqwWdSuMhUyWCNfm8x3
1vT+cag5pqRUDM9cXhGPqbtIXXHK7pfqp4LY017zWTKlz0gsgNHTwefC/e6NHGgNIyr1gAHc0KTR
noC43RbK7xMsiLMcOdrfTPz7jPth52IpDOvhi4uKUEVDh1TR3PCIfNgRYd7cqgY/dADUDkallKfE
JkrXwtEjbrXGdK2uWgqAaxKW0TyydgDlYf+AIe4tdJlEzl/FRYFmT0x4qrGznznFoMsSLetrsr8i
UY6pl09wy7fki1oyrCiW0wdLe6t/H4ubQyBOuJjp0zeSb75n2PMOYOKZHhB7NX3qwd0cMsFaiOfs
j03SpIbx6JqHUiU9k6h3WQuYKK2gcd6SKgeINsSQbDr/5iOgyD5F8143kgkDXC22N5nCQWVjgZmj
gmm/ZlIZmcELuVRA9QY40hh288yRob2FB6NV0USafRZt7Ms/lOw2JGW5JKi8Am5IIKYjY0BKzuc0
mZkU+DA65gcckOYXSWrUnTkNGe8+WrpFJrINsBiGhp6F3dnUgL0ULclUwo2A0o58VIviBr0W8QJ7
6CK/5W+CGXUEveZXW2s4Fpr/xjysh2B4vfS1p3bbMXUJgOkyK4tbtrQLCwF0pAnm6QIr0eNNWeAG
RSanCXa0qFJp0fvEHcXcuIWuSm+TOS0y5HLNEMwk8Lf9Ap6G4Cil7I1mrRWS2NcEKkU39DlIORBc
tvQGxRDXmzlNstXoXd9bhiW4lJ0ZMXXImc8knt76CSlxsUniQKcx53XZIXmKjM4rpMUSF4Ad5rVV
7W/dovLFNhOkmHU9gOgOx0Ah8rk0S8T+baDpvujCBGvWEjqvDAcHTZ//Q2c+JWNNcIAPp8Q1Ceee
ovIlAwmWlJi0wnyPleI0/tF7SjFmd7LrBNep/s/FMmLvZlaS/Z6h9ziaHUzKYAYi0GoJK5UjXJmM
ISXuG3Z6AmFBxRoGbxOfXH+KBd66LDS6ZBGeZ8hzcbNnLvdAZzfJbgiPMS9sEIyWYm3BIshYzZij
xJSCQmP/f+3KysZ6skAhHHRkXk8L/drjRAUdbsRRFxgcSeAOIDsxmiyy41TaF4uMc7vbu6Wcp99c
gIGJ/WSrRxuvyXp30bKxKq+Q8/QDNX6Nh1a1thvQzETezoUQdl3jTkGkTt4v19unEUd9re+MgDZp
EmTKbhXq0l/RjdFg6bv86Ue5qBEbBS4jhMmUxuJ0VXL9EGQ9GHhI4wfIb2CUyRXFfVefPGjygK2Q
rm1Lxz0Nd5AqceCwtra8wO94SkMlb6X2T81nsxjbqAcBZ9/Eppbc6AnaUXHTb5C45V2agIxrbyHK
+EHXsGhmPtkA6/5Iv6SEfjhG8HPAd4ssZYxznBfgrH2b4/EU3fGd+aoueF7tp2HKfMpo2KPfmBSx
NPUuXpyujc8hKvhT4rU3u2TD5pJC3hk3HoqmZO2/F5cF+c8EFRt6rYLRpYdS+8mDWqQGDhZ5mgib
gaNvlM5sF63yd+mDjVMOOWKmejEdO4PUGqRakw/TuMmVqwvvYDLqcKfLJQjs6lvPYY42aIrADTnT
h8W2LeiCzywWDhs+iZQE+mA+bzqGnQxJn1ci16LSAxd7DZEIeExWPbMh87ItiBbbuAPTg95P7SV6
c+fILYVPouNR9KLeTqzYJ0z6YDwsFmy2t8z0wMXDFJGgRyRlhCYl1q1oPeDwF3Vi/hpHEpilxEYK
+6GgfO70aFcSoAPjBiYgHIepVsCbX6NfGr/VL485d2BqQ32JwrNJxpYsXmGtDINgQFn5S3fsRvRa
CYpuUHW4cQRh0F2WtjZOsfiKkCwNp+WNktI2KxVYfEDcXZID6BMf/+/VFxmVrbEfi1FvoljkMTHZ
cFYtT63RB2sw2ErLSBONl3bE4AxxNjKV2AxFFIXET7BATepD70Znc5d3q/roDi5smt+Z6T0xIYK7
qXX5Hi0pq52+JfJuVSXJIVGHiXnop8+1Rc4hlUXFz4dZoUVLdLPenZWBQmYKaYu6fgQwjQ9dXGlQ
+pAVhIxy/EUVsa1qKpOmwjjzBzNpo1w2qBf0Z09G6hrD76kvG6Nc+wDBr/CATflebMfD8/6uQEiU
98RU/EfJE8s4mzzRtnUiPE6p2r7nBf7SbXMaHoF4AyoxKpWI2/3upl60FVxkGVyjpa7YKjKGlZe/
tjN6D/kERPBAlArL/NQdvnRLitCd9z6YMLgSuVOivy17fCnHdlKbPf/lOJ2aNaqOQvPAI/UU7x/S
Hb2/5UWozP1+3EvkS1deTmycJ5pP5x0XMXK3TQZqO9UdE4ign6LledVU8VjldKY2220khX1QgmPW
E9gCJSYypwH55vKqr53q/p4jSHEDyo/fWgz3Y7iNmIy8lHD9YmtQ3/HZVn00I4vJA6Kn4YNVPPxu
g4XC1i73ljvUOLvJ3a8xZnD0jQdvGA1YNW4Nq7myVWkdRvq2u1FWh2ZLQu0edhx6J4OzyMdjTpcN
bkoVD4Cakuex1k773u2Ga4BzPI/Fwdcy7/eeZvcENeuBEEzBNMdY37fSjI6JsRS2BTUG1/V3IxaQ
mes7KLFuyBSXzIs/mV/MBB0/CeAjC3R7ydiaMHd3eH2JGh1D+jGLsoaQ/BP5hiyezJgmpQqUKdg2
HBHwQP0ednAuaZ2S2/Rox1Opu0O25zJvvTIetDKYvcQdzCL8URo7aCD5MfC1R46CdmkKpEo1XCup
p1Ml0tysg1Ft4Tq+d0ZzfEZVY5Ivk2AQWKZVQMZ+EXQW3gvav8YHQer3Q9Bcs1ohNDOGtYNKI1tc
7edXP+2zJrwZNn4sN/55Rp+eCn+w2km9nBF+/SYFj4LLGqrA3MaM9HS6+bsrNuAnXbJOrAvC6HsN
mBPdZ3paeLIjNZPjdo4q2+37Z0A+3ijj4Qmhzoe6hVBZFvw0s3Kc5Oz5dzrw/96OTGEBXibm6ZMH
kT2N0nwnW/2UVmzY/+jIgSsQJwa2rLPc3TLLygh1M/PYPnKPEc44p7YuPf0bhjJI7UYFQcPE9CRW
//T3C9u4B2DmhNPgnMD4XJvmhumlhI0JYBeFqCqN9wgaSvpnakBmrlqYCiEgt3hcEzMXmVKWpzYt
1wMO6JdQiplKyo5ygKT6/r3T8O+JXWZtdHCeBDBGHRQOBGoZgMRCHKcAUdaMeSKZ0AWiNjfbcmRJ
vxm2dcpFXg87EGjhjjKYnDJpJcU4wdmegvmeDWKEthGSXxwn7VHlyA7iOoPEqD9bWPkIBIBH4hcj
8UlZrYU4nweqyRvugeGRMDZWRSaz96hn9788vxSbwmVQYcFYOQaVow3tDK0KAljA8/RX10Sq+Qev
FVPrhYTZwyA+JNHJHIqepfNE4Ip9VlgWwQdepVdpnB9biMbnRhXzxtMa6KKq0nV40Sv0stiQLQSF
50J/dJq6cUUf+50ZUqC4tVZtrFt+hEumovu1bR8TObkpVUEgCtcvYPPnOzSchGgG6shvqoIkj14e
xJ3SAHE3GqSjOYxpUIQOWNf9qiEe7KnkpofM7KkohX4PLklS3V8DeJTOCKRnd/2jIE38vWZ/AjZ2
FFzrLm0/xG+SazGgYIohshBHxLIMeJ3a7lqw0rN+p2lo58nhvC8R8uDDhQU+OyhIf5BmLg7Bva/t
m8S328U3J4V9fXphXH5W9Hhu0wYDfm3VJXoKod8zbEpA+1MLhGgIoEPq+ku04RMNYKguGvmDUDrL
1xXe3a6WwkvoLwf/4NtP1tmxVQNP5Lmi4FivpPDAVTMffOP6BCW+lAuiBYjL4sLqb5Cgj6NFQ8Cr
caJzspaXWue0i7tkMSU9jE4dyz1msCYo66fELkTiSuN1uoOcmbP0WAHzla2UJExOZA4xG+ww172s
fUzwigh91eowYkuWrLiOP4scNHgZhWB7V7Sm0hkIsjDXY+v4c06ISVNkUJsJq4zaHtYpqQeKTHO/
OquKVjuSosZUOnNLXVbzX2RSNV302dQmkYcy2nuyopyMgubGitGMECKeF8GP4t/HgEYSyZGfR2Q/
43ZbyrwqCUy93PR/J9kg3q9Za0SuV/xq68ecbrK82mHnKwZO6Ld1PD4J/l1zIIS3F02XSOq8VSRO
x1r5i3h6lyvmQUdt2osRmMT11qOmVJMk4TQ1NUOyvOglfR0T703XktP1mdOIL1d6ZUJ4bXo6iN1+
yKe/pQKaOQn2/mcBGk9Y31NK1CvW2srBWHwf3AChCQ0mNT1IsnZx4+2BzvDCwaJZOCku5UYfNucY
62L2+WVQCfv0eT6GNW5MxbG8XflM42TDRhD09Nk2jR/neQMWwrXVGzJu68FybuX5Afg2A+1uOLUz
JFZSZIZKNJ5OgKeZsIK/aHc7ay2iABtOu+22J5C6ZNOLktj/1QDdTgrxurdVIxxYfQHvtfcP7N4m
BADGHjU2qXvWXK54QC8c890BOjkLpsji0T73xLOXbLH/W92FwnyzFbCof5iT7WeVEGRk+96a7jUc
IP3VHylQof9Og6WcOV5I9bE6NeBkJIcp8G9Ds4GlQnzA1PrOoA6MzsFtJ1FBUqGOASE6QSBc/1fN
/YgCZyx/td1w9g2BU2tTWksWV67YzvfPb2LxJ4ZMaeFTM12PA6/+uvbHhW03v5sIEU+nV6OjAYmh
1ov4b8+AlcPn4QQZzxHjQlDGoMkUYm2+iXn9+DU3AfOcO4+uBAH5K9d2ySPqJjtW+ejnm3O5QU2S
zc4AZv4zZqecG0776UH/mVInRBDfuaYpDg+6sJwqBruJzCcp7+8YIWNVbfLI7IyskvyKYxui1ymq
1CwZ2+dlheDPaXC/cLUOwovpPaqmymBdghWlKAYbObiAOjUTr+O2bkq1Eaz1DN3jj+eM7pC8ndx5
/cjnaTBYENwIN5rswckAkyanmRIUNAswdxukrYhNuVe7EBPgAmLoMbGSUUmJ3w1Cim7HSgNUOgfI
fW6wpSr90HqoaGmQuinHAYDhBFx0MAj1SBJx/Xv+vJaqdCA4gholVsGp9NEG+XHWCZ4ytm8gcm/y
UgLA6Iym2Ak3/6Su4J7i9AkKr4pXRo/irH+HQpxUs68gfm8B9NJRcvHzCi6MkImPyNw9aJsz/l+H
cuNscAT/CcdeXhZsnDxod1hPslkr5sG0fd/vTk1+2147T69K5zrmaXQQWNGCLCLyUasBDgfL68p1
gFfQijnH3DloIPuKmlgnD/rbJnYCmHKeTAAWe87tVQnGb+z9JnbGJprTeZ5Ro2UAaDbpnx+BHNpX
GVvnf0MLghkPH8cJsWOyoeHhlLqiX+qznucUvSgTpENpNbqofULxYlStRv/2vvdPqSajipj+tS2S
iEKPv0fhKzGRi/NlVzGpun/XYPAu1cwBUrmkMayuxgy9T97uJ7oXNKNtXbL7ra8nE9rE0O60A4+b
J4TdLrYU2XQm+xabzpX0c2sKSlph1NYQqpMW6cigJJzqCgxubS4K37PaufBCytMeEt5s7/HUKGcs
fpHD/tmlOrvOPkvxOSU/mctXGjFPRSpwEPZhHUnPxFysSFIqM4gzGER7G9i4hVENcqDEGA3U9ice
nWQ+9TGam/t4XpO//zABaWorrZXKvMi+9Th31Ed/TzCGCkQ/rBZR8D2KYby1WrttqtSQQxRytm+n
5zN0qkF+hw0tqifyjv2ElmohKgFTHpJjMjhXxQKcB+RGz9FHZcEloxrNXtwD1RHaKgfzm/yGbg+S
j3C1PSzj6bFit06pw0opYpij3C4qm/2OPw2uVaFLyEvJ8hw8WFkv+YP6Sh7ZYCTxbfYq1UU3PG21
o1SyzBP4jexcicIbRkLJtyqxFNXQ5wQDybOXyFHn/65CUd0IzNHJDfrSxAUU/rBl7aaaO3kAOccm
zIR/0XvaEnsKwRPlo6u9dH/XrolgiKQesRqz6rBGd1vKCVjHg1n8gFRDm1jiqGM3ldoMc4e4aawx
LyHP1s05gbXtJkVkh2xuyVTYuZMt/vcwuJ3EjASqqkzHH/oMd2Dh2ZeWDY/60/EtWf8mBE4xTSMT
VLcQD9ZWTas9GeCtB24frNSmStAbINRxnqbJbxtK/VCbJkh716bTlKKQQEvDN1r8CBsp8pG3K/H8
Jv7pwcVGxilgNLcvSzubgx5KCFhfxxJpgrtn4Tgu/107FauF/i7whumvNKHpDPUCZUNXXvHujGyK
Sq5lHhUlMlrbk8h5c+ya++azIgHAFwSPPKdkWLzuQRsJ4e/cTEEInORUVq9Cozn6Ck9qFzHGVWHc
51l1ue0lKOoKnfnMPYN+pxbLNOKSWnCIEvbX/jNNaGpKcMTiIBS86/VdiKyrN4I4HpqBuSlHWWDK
EhktO4VMLZqP+PzIbLPCDjVLI3yn9lCNsc7zTEL7SYrJuPCRKA82Ke/IoCGQtbv0N9reRmt6ao9h
Pex3FkXgxWkgwTBgZDA5Oklxgsn+I5aE1KnZeppaOAK/fRyWHbGj9VnEzzhPhFQ+4p7unV0jrkRP
cGFes1hRCBRMoWnBxLcng1XvhMx51E46866dEz5o/P3chY/Wy9nQaw5mI7mPEu9GcOA1f5JXDzjm
6Bd2vtmJb5R8Cdbp+p4KN2E7IT16vSKAc7jOOlzHUpGF7kVXJPo+vUsY0r2wlibRNxx/On182l63
1Gs1QFLMwXZuk/eW+N0lr+efnQP7RqkbjmatJfd5aAP5XDNMgR9qXuIRD/2IEt8rhrZJOjFyGKdg
+GqVjlN5wXTMqW3vi0XAYIEbAZgSOnWfSjAjStMYOIKP+xH70sk6YDPRu/NmxUF9OUdR8sG7UDJr
oCMNQzhpeOj5YU3WbJtMfW3vm5S62V7lwFCQ8R5iA/LTMHsDWAW7v8lrrOodooCHdclAJlyWb5Ig
d5v3vsk7Grbg/MnNVdSztgIElnEBKIGukC9pFZSN8GOUe2H7vPH2simOI/WFUPEkGqbWHhLbdr/M
LWuM1A9Y6qAwRSEOR+wQ0uWlsS2p8+ap32VUhsQouYDFTpsi3l5lHoTAfyMd241yXTKa5XZmscOu
UOqXD+qK7pLd2tWzJiYrvqyHR5X8sVCRZUr3XHljjcFriLzRl4ea/brctq29W/EvDwGDpQPG6ggc
eOLFSdPl0M+eKO5e+1fTVR0oBgqUu5QXQE04f6GWpDIYqXZDhiLJ1MlN1nzqWEDBivt8MA6Oqu3+
VlEQuBmXftDuJObfMIMeTeiyB6pSdeIyo9C1pmBakTGpgM7n9vSytC8FWKBod+gGyPPE4XSB13Z3
YwFDBLCvPSWTS1rGGg5OMIFP1RYFbFzcyX5SUF1Ye5Wk5hchvIbvZge0yHF90EbaskHSmOyUc+d5
6N4z35v52t9KItF1ZBbDySHB7NIpKYLaEr/Ghl36/FTEbmfx16x8H0llzGZqyteqQPFfO53EICzo
TS5tZng9WB1G1rTCaJUZ9JXA/zLpDQHbrzfAPrRq6VUndemUuusewqyjQdKUdz16W6nGF13phDHu
ax5xa5mE0xRh/7Lt8oA7wYea0iDUn/itFKfvW0TYSjo8pypqBVBdFwovpuLxgylbti5x3wWaBMta
iFS0IUtBeEF8H2BHVfuG4iZYDx/oguwBDBvYyFEaSNyhy8vw82jmELGR+7vL7pgxEUibbVI7VAYF
BylBmWTAE3CUV0b8anNj6p7+gIw7p0hLuaoAT7z4AO6neLaO98hJOm7XnidGSYL5ef6o5J+vW5oy
LgLSu0uU8deML6vGu13LySiW8ncaCzBwm3uZUzKThrxQ/Ez6OpJCou120YdYBx2OWYxxYVX9tGft
QpnZLGkgta0OmGdLM0wJkJjwfAN2N1Hp+XPBUa60KjypwnYi6wQPJWcUifisRnmoR4+8hKZ1ysJ4
4/dpDRMWTtBMSX1EXka/4jVtSdwotcJMwezqB9ymlCmM3r92ETdBMXeX0QS2H9ORB3AOOJykPX4F
La33zA9N5AvzP0F8pMi+3zg/sacS/sKePzwmmnHW8Tfg3cew0SjoagQCZnpVwppkNoI92OOky2WJ
AAWsx05VUXZNiJn5gQD3iY70ztreCNY5bpp7LxbQbvYSmJGMhY8ftQo+S/j8vgvCF5bFlpSWQl7e
FIgTqCg6JqrctkWonaFl3I7OYpJ0lX/whSDi/spWPDQ4yEXr24b4qV8c9c0ERO1AC0wfTQ/chjOs
O1mnUtttto/BZOafXUecWULg5UobRvYotZtPrPWZanoWgOHZyVokaAc6SqgiKLtrvTmTPs73eosN
6zR20Wywr18FUTj4xS6qrFb5FDWq9avE3dB5XmrhHyxCQba50cAdWh9tLiD0SvZOsmERC/u21A6E
a0T0YGnvYlOKsYl7W0wVVqkRUr4JxmXXcq0/n4F3IvS1mcSzu19DcFmOk9YdDWP3/nxf3bfN8HqU
EpVXddfsXQ/N832etR0GcpejAv/U/vIk8RN5vDiSyZRIevK6pVOwYYZZ7nt3weyf3LpPi5uMcHIi
iqH1gZvl8UU6PDljnSWkCSeZyQDcDADuAN3n0WcuPhv+AIUJrXr5DeQnbC/75w6pBoqlkiZwKnRs
dXyMrYJvXJmUIIEbXl4N29MOyIfk0wE8Sya//0JPLVFKpfMUtP6O3zQv+3QYJm78nsAMJQvQ9ZV1
fcEmaRMrtYKI8imiqq+UdCdToOvBnO4jymWk8PfjEs0RoXMUvxpz8ASM9iwQshW0QjU7EI0X/3gE
a4vZeLIYT9xCZMxdyS1ggLIo6hqj9RxM4NQSBAOCZC9DGc3XIJKClxyPsE3SPuHEmbq0iQDuc76Q
jdyXuKxfMY95duLOSzPHvVJemciqQc2rddreqPl7ezIkoHWP/QMImfntH4J8nHdtCOUkbP0kKBhu
oHvAc7vFt6ZDdQ20mvc2UkVMu2gE0GrNiD45t1KbB5A187ByzPblDEJz5k7zDoWa38Ub5F3Z+amf
xWODMXqcIz/eyjaEHgq5EAc2W04tKDlPiMFk0LHqn7CE/qwis/FN64JzDQVXqeAKGjKPixws/9kQ
QklTwAzC9YlX0ZKtw0tKzfRCmhF5Y3ngq5sj7b0mRnBxRVkqA3yfBiJyPT0c1i/poWMJA1AQZX58
HS00VWKDfovat2hNXIcDiJdm7wMJIo+XFZCAwotPauKxpUv1B5kW5XFQdqIgRxooUrAAOO7k7Zij
36vIUULGB/OlTZ5Uj9GqcXB1h/5rLXWWRPVeMBKK/9e4KDzYoTwzjws+HfHGlo2Reakhv2GcHnGS
RnItj+jUKP9NUa2A30+HLqHG6771TgFkhX+d+8phZv5oVULIDDm6//8Wf6sbTEHCQ+QSVtFZZgag
OTVBkCsBBkU5SDzysRBsFHwAMu5Kg1XSswvsCqPeJ9FgVKXr78sdl5GeR6oF/EAYrbD86wXXOc2h
zdeGDQk6tCI5RnjcHypzdflrHbqr02BNoyibX/WhUj6c7yxII4xM+2YIlKMJjplBrGTf3n2O9CIP
g28h9+kjJNUzjAMa0cY4zDmWu9B4aOGWsbpad0TTmnldvSkfhEo8p8IyLu5ka1iyv13BWqq9K6XF
PFzB0gTi3XcP3taqFshAONhZu5jKyY7fcy7iJ+MezvEKJ3CfivskKThFDC9402StIlPhjk65Mw0q
rCV+8H7Zd6gCgdbukXfPQ5m0rzUgCEPDBLEhOAPx8d6CYBa8HArL930TvhPqr40mPIiPpcJCZc3t
GiWA5YMNWvs1CerWMx2m9kzRKVaqJR1NoW0eg9iRUXSCIaluFx0LCF81hbOSfh+LaiYhbusKwq0P
Yg3wduPbybVFnfmTGPtMlhznP3bsyQSAFj+ns96PCRxU+r/JZb6iZUhD6E7boKvX4jYqxGG3dMEr
Z+drUSCffc5ep8lMEVXtK0OLReNZnRmqik2bUq628ewEUglIW4orZR94QUR3C0ReenIMdNyX/FMu
StJSnOgx6XSKiUiqyF4w3i6rTfRxSQAe0zJRJR60IyS6DFu2BucvtKKuRZYTFAbT0H9K95ExabNb
zRUoSo8YzBpAiRSdUUp3pO3n0ePTrgZDyyTyJKe0iP8+4A9vWolaK8LRQeuko+GHkaLivZx6V7cR
sUDkc0kqragKLaxJftLi2bReybysoUx64AZirp9jjd5D43LRQzsyEg5mlrkxVp2DD75JeIrX69je
HoVqLhELx+ZuHu996crsKHzl2gPBrrShE1ZGKJHiLq8+UomB0ZLuEQXoLoVD2niwwkUEEMH88p9b
kgdKsp20314WbKjegx2v2Jes1nxWDNptVNEBPgtwvCZXcKVKojzoQaEKj1P2qZ9cs5n2LBXKF7il
zYRqGhgAUeCwNikx+KlMschknzOaKKxuoGDpwjVKdgCXVH9CsU+rf1+RfwqHXepS/oPZZBWsa3QT
o1M8AbVfGM1NMpSsyFhwwzcgHPfbY8Z6i5G2RILsNDMmyPX6DXHUkDUG19OrQzgCnc6Fc488p6ja
lKDYSZ/5hBjLDu8MA1Xm/sr5mX8TyVH52C5xZZKfML+baSu4pByv5aOYvy46JpdyzCAeN6CqbI66
PQ5Vj3vDdvpmOHah56mEbiaBSgdy21uo/Qe+h8WCcPmiiZ7CIubGtUVhrl/PKJpIa1MAqkRjoy/d
VfWreJW/fNvGBv+Q/lLo/vCctGcPk6D33DuNFNpuTagGXy0QYx0rrMfumVW4ddkIKNXk2ZAqOYa/
4RvS9Qse2MNPnoWik0tE2qDzYDK/k3AkJaMKlaioaGj92BYm1aKKDT6keceDTVsv71ThWaKcOqAG
KlGf8LhaRjeQC6wpudJovBNiCouzPah3A4LrPjtplLd2AvenrC/Optv548GT/WSx0fwzBrMjY11p
shLEv1Nf5HO01IxVRJmo24kjqSStrV4L5zIb2Hla5C4DpkUF2/wOYnnNcDG8QCuldGvBGruVwvih
d+6RrGZtZJJ47GXz0FwvH0UOoOovjOYTPEwBlACYXhOwl42kBFSDbx/Wpb6u5F7g0zWFppYZb19w
w2Hzdd7WKvxpJtO0WiUaIdr7eAbCx48u6FE3fv07+WiKQeazYXOL1ZICKgPEFtbttjRfHluPaaKA
n9XHnCiUMHXZO5gQFzqvSHPMedy2k+uWaT6Ilg0ty9pqtrTItmdnTKWmKXsBriOeZiPlwsTBqY63
Vy1LyGRIo+fb6XjWEszV2g3OYVBQwx3M5/+nJoj6zNaEFpwjmmseY20q0q0iaByEp3O99GqmdN2u
OMZL7Cklc/05Bj/dEKrsVEUfYZUsSfvq0S9E8E1CXHFbH+RfJ/zd23UQzRsuMNlVDBYbcNtU1CdI
e8YtO54vNzrPR6O72MjiftCvL9wrnegZSgSnvjewFmnQwYn8G6acs4/WI6uH4oIboE3vBYXiV8Mz
fQhQmGoSnxyTKsji8NOXFvyAKDX2OcUUKJ9V1bd+NGf1u9GZVIULDmhDV/su48uKEJljUSMl6LYp
8BnrGBJPYwMtiI198ih3c1O/+IdcxVdu1TH1KgQQSdORvsnmI29u2BNc1mTIvlLNwPRPHBG69kcV
48egKJKby019wKNSRKK9vPJKvH36I3hGnvekWca4zToRuXsy0SgWRfHZs/bT40C3BtYk9NAk9tJ2
8qNIAI37MCUA4mzkXSyfd9o6f/KoC435+n3BjG59z1uf7dd9C9nUJGl1nXNLA4fNZZzvRFyQ++gi
jZoDZntIqA6r4/RdG4Oa2tnId14/zEf75G1WKzDq3mT6BWfp6OPArf76uniE4efkxB+Seq87xsiM
BHl5k8mZD2PqeBUoXqUX0/i9G0ht+Dd3r13KWLKKnZ1Z4NlzkC/SotjtJiQxXDZSe1cQ/v6EPYnk
YfsydpjHLyKl2VI0edV58v4C2KoC4ORKETP/nBhW9OeMVDvH9/t8PA4f2NUMjEzGWQcz+i31cY3u
hjoG599W8b+HePmiyMJsIh80dlY747G3GSYAF0AxsiM3hPpQBOe/SSFLa4ovB3TaupQXwLVMYXK3
jJy1D9s85BB8idcerTRurNxuEBz4dakwJBJYK+4m0cKIHiqS2KzSmQ53AgOE6RpwZ7ADq7Bm8Jbr
hH4cwtK2446Z8Vc8jAR08ee9Ux4qyCfvPJnP3x69FgzqEQKL9+S+2rIiii+D11OFuWp8KPUdrSzt
Qe8xzjcD2pzRwL/zFQsRGI38dLiSui2nA0UXtbqykCYCUHbcFKw5yWyirWYLzrQZDffHzMq115gZ
stJp0ModhE7WLGoGsLxMHJV5HXMs5naJQz4x1W+PsLH8bJEtcIJya0bG/bQaYznt0T9TZ0Cang3D
JfZuUCSg5lGhZg/tVh9477n/fT41E2U0hZBX3O9WqFTQdkkjUCXUWqo9Dg1Na2Jf2MbRSVEJDByN
nZ0M4Ru4LQzsejswxc6Z60WEqj/6tSA3JxBFd/9rty4/9lj5xl2QvZSP/T5fgtqW8ddxwFk6Xm70
GJe1d6gZqWhXqb1/GfQQMShHTyuOXvBP0cLKKDNk8ICv+YYby2FP9yScvGdnGMklzTKpFQNCqrR9
qA+kpkW5Y+32jZfSZ1Qojd09okc5pbFrwFd4SW1tWb/I/rOg3bP4leWOvJz4wePxgPjsKpMsEvGt
UgdCylya/QL2knwM1AyGUo7EM0DN3Vf3cI1MPq6CgCF32wcrIzrRIfijuUheF4VKffg24YOE/McV
aYJ68ebaAr5UPkVCorTswKcuD27J1yZ3M5d+w6Rp63YYX+9qiVFC/nZzU33J3dDcPsl3Mv4KeuY5
LpHTALi4bcEetvgT6ozO3Ma7topXM4nqFUXusJ9CjaNpp80ZrW5eDPyjH4q1+po1tOTt27N+mNq9
5zdyQTwoULvW7NWKAqoQrfnh8RuG4QVvcmdBFR7wlkgZ8S3ipeNhKvhqlcU3AX0QUFCp/q2qMrRa
dMCn+Bx7e7cFJ7K18ymhY1x9eTCZRf+yICAGyo5fN1zX27i3/W/Ks37p0Lffdq3s85sG6xlpbT+4
gDL0a5RjHCKdSdfX50SxQD1IEJ2qUJQ3aGaKmf74kQctPQbUvKTm04Wge7neqOfR0ZJYAp3hm1nU
nEJZvf/XXnAOvDZJx1zM1TDDnuOfkrZyjmtiDvqK7TsXDC6fANQRswS/qTCTxlNfb25feza/cYKp
Ou+vAA52ALMsd2guv/6rDt+LKs9S2zhScQ90xmomzdFyFWpoZNRSGVRXSdJRSgJqeCOedRbCtM3t
fJMEs2FkDb6u2qMmYt9DD3OUuq+Uf3X5CtwpDD5HfC3mW8h5pqs6/WkJhuY4YEPmglGTxXBdU5KY
1dJzLSwdkjS/yHL05wmvCK4NyfHZEFy6fq0recdcgE3XDfDPMgLnkQNPsZGJ4xWgiAthdU1/P/bF
j+xh3RX57Qa6sBJik7K1z08YO2Br2wn1PIkZ2I6JIlC6c3CPMgjUS/bqElGV8UF9MtwZX8Emj8Dj
UzuBTbE2JcOyCw76gsW1CF4hneoQnFn77X1JRjs0hF/lG6edh1J/Nl3f2A1CYa8aZLDq3pUFQUhR
1AJCyX32QA0FhubSd8qLuOLrA0tFf6rT4+ismp0h87+QZjR9zDwXugVryskRYM4L8FQO6cBkPNw1
On66ikUhXo738sbOXmDPwMPo5fAgxgqS2+lzbhPhlyspyo39T6UMQxsxFvxlOlWDg0wvaRidydoC
1hUtCkBJwfXN0tGR/V7m9t3Omis2Xnm71RIFxQ0Co+YzhT1tpWm6ugn0KmYR3pxcrrHXr8cQUm+h
2tbOW5ipAeS3DM8PLAehV9Eilldge6l2r9DE3FSoq9C7M4pIvLaj26kojkHkeD7gL2Q+3bNF9aog
W8U4ZA3OKsrw5e5joue33CDAOpuu0pxo1jwMBLBODPq267WUcAjVumeAEHFSnjtiOxmV5VkUvkuk
LtrV+IVy2Gdz1hGLx1JSwlXFYcuPbmHz9qWPHGdMJiK9sOcsYeexHD0xmwCkHf0EFuw+WWJWHOtt
fqR2WFylrvPp/s7isje6OscE8b4G5WjW7gxkV7v0bblX5Waefne8JXFiTQTA6ZRWmzkfHcr7Esj/
tGkvOwGQPdFVnV0HKUXhbWv47xUNNBhZNUrxDmZ0j9V1E4iQkQwwLUrYOYgpwP5yT7n+9yOc6H8/
tAaH9L07mut3wSa27d+Q/Y2EQOQSqVdp7jzaxO2G2k2qGGkP6XWlc0R7tnKqwbTqeWrqvAvd/SSX
Pb/gv/vptepA22xZgF4GwfahXD36LaYPq14OmgQjRoftHrx9Dj6o+FLedytg4cQRGz3w7Oz7JYxM
rw3Wf+3BoDcNtQ9hOT+gLggo4KjGgPLwFOTB7G4QsXbsKn5b2ISoxsd7bfwBbA5WAMI5DV6F0/W4
WVfLmu9+tnQswk7t2/ccRXAOVJtYztnLq1LFY0J0KO8nGJQK+i8nTcBrWwbJos39a3R0+3Opgete
YcbGsNLkIb+3AtY4+5xrSPttAPaPga0LRRqjDahuGjcovMC//47IseQ/Op1IaA+f4CuQlHVggVKY
JlhzOuNyHbeCeKZXt7K9Vz5oJ0jG898jwThTR2ndYIUTzaJGsKicyE4c7lDF5zCT0sLJ4nYi47ex
zenlK1Kd/JxYb70BO3UAE4ZZ5sArQHhVkdquEpwNe1ExFreXx02UTxbGiLn7i071NA3WlI78LDq4
QVjagxcqAeigpWfdzNcJC7z3D3JsaJsUOVvqXG0NzU71v0Q0eRC65xzcjRv+SjVOJuqsOzqUnV3S
5Bs2/lA9uh2a0tmWUDU646hcs7GDS/6PFvx3taakIj2ZJMQ+EfhzcUeVuM/cVxkVQXLNxaXPF++g
oJEn2cElTJSOYSYA6hbFfVyeo1znDkkS9stEQU7nNLYA6XweLqHPyRRJ8nRt1qk/7fk3RPJRbE+N
6A4oLogcxNmfJOZnwFpWLDu1WiPdF9XsRdGpsd/ydiWSZJuzQU1aALh8KKxFra6QXJ5xikP1oT6s
1rSMWjoEkX8c5bl907hb4JKxT5DwSEbEBemLzYgF2sgJ/6uJuTof/mXlkij2w0FN50VSP5mGuZRc
RiJ+X8HzqmIsyS9caxHVThgH0kJKBZaC648PJUlh0GfG1o41/kV1gNHPZ0ktcvxsoOPFnKQ5Onyl
6vo95xUGrpMTPJhZNNE3X0Om8FCnaPmWW4eWb3KyhEzxsso2j9wtA9XXADKvSgYCpgObxppoW3XI
YlA62aPkX2Cal0B/ekEBMqa/AVKC8t0E9OavOj6Xqtng7dGezBo6AwVNZ2doCcoQsWR3yfLknnWk
k9Rz/MdPdwfxZE4+bcrKt/zh0gkJkjd3nVePPEfirkgk/yPXqWWzvR6ALDsO8hdk1JiSCwk8r3B0
Cl5fGV3L/iTLuw2D4sAG+Wwddf7t+FQngwtmdQ4TazvRancQQJazz91MXvRsWGetf2KEijQabGnC
p4P4N1q8IrOBZm+rE3xvkPP9wuXwNTmKWHcCQ6j8LZ4xgb0rp1VH2B/7CSLmEbeDKu7e10xj9qpn
DQl+iHdkrjRNb/tbj13hxfHu9UDP8wZZg2cZ9BZiHI409vKId+GGRu9gbmjo8TFxg/rWhplLFpvp
ICFH/KKRk4tuP3kvEzriGv8hKtf38ksjXpdVtWZRzpuw6zeWL0AEkpI7tW0Uuorz5W9mOHLmj8d8
VA3cYkFv10pe81zGBFY5f+RUa1iYg1VRSi5ZIQGaO+frI5HNKJIDaYGHmLBgE+F/sNm0yjknNcBP
/1G8GvSNF7tOdAAw0K0czzXzvVqrCLalXYl1/zqlzBQj5m9eECVeQfd2sAFUuDS5HxQ6Ib5MsLyt
C9VYKZ3xnBmBowOcnwDurnmSmB1LN7gFmRkyHxkaz80PXHxse10ip7E5eNLck1QH8tJbqfb0WYtR
11TjG6NqVGMtGr+9GzVyWYjrEE/uHBWyr3Ls7xTEkcqwY2fgV62kX4/ISdvJDZ2JUVucPj8/2pYz
/ULy4E/g5mPtD+/MA4qZ/GhB82REdvUHXF70lrRWuN2hhfGOltNvcChUyor+xQOAoWRD5X/CyFvA
o31YR+Gqxhbhh1+3k4vkNw/8ElCdQXZsCjKXpaiy8MbZQ9Ovuhp8/cGeFSpozuCdi8fVqYLYvpjD
ydzKodvSPS/ESfRnmw0DnyoWke/ErDerDMgtGtvnhOmo7+T0e5w6LW1K0ManBAspma9/9aiPXQSF
V9iURqI7B1QhGHSHpfiw6YP3tE7ST6EyJaXu8KnS0GVAECQRkgAoV+2hapzNC0fmLfX8nzLAjeKQ
+AZ2RFzuc9td+Yh8SK1WUScet458PJVXAyHdanIe8vq+2NCApCNYyZu+zVFH4OCzfWRcwavR8+CU
e1eKWd2hyM92dOlwqnGr7fqq2AQcaUlnCk99bh6hkchG3mF4brG8fTR7XmCHy9LvAqxQTSY/z1zY
cLRjG0gCROyp0wTDgkri8+eN6+XWoRXuml57tTCTO8gLd/pnkED+7PNTpFIB3Dm9TwIiBm5Cj+SE
eNN6elHqLbaSF1FcjzEjZ6nGdpeKN6rYHaVrCWqgkzqyAsCJzMZtEPrhMUo3apb1hslQv9tvFF64
KmyjetibLjdNHUz6zuVdUGO7PHHKOcxOaefqm8xG1CkyeFQSQEVyt8X+y4bgQjNSmoRfJIhfjGwe
5p/yWbsq5BEMCP7ljMN3OPEN/+sUGt6SYJJbvru/2y/n5YfwUPkaSX+f19H8jN93qiPaeJnVjATt
hiCVxwdVn5Jw+ACJddDcS3wdSGe+DdZo79+pqLxG+/9/tTpRGGdEM7V3BZ1G3r6Xt2wOCZ7BRgCC
ML+gCHwIoxewABEx0uq0VHiML+5dYYFRh9Z2pJjgBUVbOuBfVwE/FjgdjokdJeMhH0ahGjG+tFwy
WxwiV7CvKlPnsJbdrr86M5QE3q6mSGWfVP0qsNVWQc6DhnLV3w+kJQUMrDvBQV0geLzOpB7702bW
KWa55RgFGEKgr89vXBX+7FhsGwBZoh8Hli6AE6UD/UNE9I4zf5VlSbS50q62RLRFblIdcdNwt3CR
aMnNLSbPdS+edK+qtCgSqmyNbhx/vDMBA7RkepwURfdY/pfj1ZoeuFsWOEKso9qjzsHWoyyu7nl3
yX+OWfBZ4MVbPTxYC4+ChbAMq5yc/bqaLEHmH6qG1SCLKmfWRE1okW2HWNVq6pLcV9EnePGzedvQ
yDtlnMNoDWvzjPoOBhQOKkMiqN1ndL2vs5Q9rJm6P9Mt94q85Dih7yDDJTP74heYOUJy6RTuo4kP
KCHGabAoTeP8evatTRMGuYyLYs8HcWIuO59bx4E9w2a5d9/9wYVNCJmoKMu710UGn2FLb1MVmNUK
UAmnvSlteTKvonSjHWDRzrNcAm2ILCYzzAfEu2mhWT9APU7L1pAEZ1gkiW7X9GRWtsIY430HIFCT
2diAdIH7KYd1HLFe4TE8JA6rx5FGK+gfzEXn3fkaEoH1kbVwmPyPZ7A7nhR8353QdV/uxq950iTL
TtZvJUkT2KBh7oOHLsBYS9wPvrlyenDK64WfvpBliA1BW8sVulGztXMTU6KhRv7HstKyqs+mGgPs
yQzrZ+j6GiLcsP8FqWO2iZSzvORV88aAizpLqfMEaAtp+qrD7cfEC/wgjfPpYPoYJVrLGcczT71s
m7Or/Rpp4ayUVQZ0Kwkm1CPV4ch2F83zJTb1zV8vOZ852YmweMp7ppY2I0Z+jL8jU2iTVIwuVmD5
DujcAGb6wVBy9fNZ5tgQuR3w0UEcO+ikqyITq5PENC/Ru6jkq9Gd9xvDz+PViBCpVau0xpcIV7z+
4lGkdlzXyQwvy5pca1rzLxx1M9iOMOXwo41Hvt75FSbJKE/7rKgtwFcbK7FqzfEltmFGo9/35sAI
NDqLtFUlQ58wpAHeqeslsYmTu3S28C+0fHHocX1bLt/e87KJycU8N6Lqex1Hv16FWF5ECctQBI3V
VRyGsrp8sJqYNm/jUyJJDDNKUCXGLYGNy3YLoKDeNUnvLr139m2WIAE76ANd6k0Rv6AIAQs0Cdro
wGUUgLiAou0UZ0G5g3ZjdIZd61/iSm8adK1ERqbppp1rB7zGfPqxLQh9MiEdcUPKECAP3hTWlLhl
rBZUcskqdunA3b+vfM+gjSip9m/ve7++IgZoD52nEIhR8bLV7GAN3cowCwkYOOnTaSJVlYticOXJ
KYVdLBywS/JGhMiSqvzD6od5PJFaeHYkQVR/RY3ZAhQWD8lYjsqbhtuuPmkGYo2bj5779gCStZce
3T9fmUerChPGP6YHHRwm5VICHUokfCu0ZQbZQSasCts/NosQ3jzxxBZsWvCtH8HwZ+PhXWXMoKVE
E0g+kWgG5Kts482Nrsp8uLhK/NyHUVgeZzmZ9uiompjQlXk55APOjmba48Ot+QgEE2szHJyInUex
n0kKonttARDWyROwD+m7OKtH8R3HheN6B2oaI2J99CejqwLpAn2Sb8Q3Pr36tWE44WFRPLMsZWWM
cy/aErddF4Ptouyy8fPQomXN7gQa9ArIY2jVpxvqz0BwfXRfJ0s3bYAl84zEvm+NcFAdvV0fMRFi
pyg9ycxrLkiau5Quh/zYAXZXD/J/DY+cD+FkihiJJvzBo8d7zTgAW1S/n5dQ5osmFcbZ/epXILLN
ltpWVTgEUKVhFPaW7acwPYu99/IZFaQpV/UTOk5xzWrp9lLTUo+4r67lsvvApZGf2UUgG556bVQq
E0Vdz/4uV17FkoyJ/1ycYKnpfQj0WlGT0/0z2gLyadyhz2MyynemSYHKG3q3u3gvMUf9N2AP1qpZ
yqpfbcvRtIijNPjL6Nb5YnMwkM2E36WNikaIsRu6nS12zg2Nrj2kNT53K5ex7sKUUDnud6QaV0s5
8wtIZFrlWmYYDclc3KHqi5Z0YOG6+eNwyH4owqUm0mjHkNjFVHrH6HWuTRfc22DaLrtgeyhmtKI3
2nJsUWsYSDg+I3uuWHFGc1C3lRMVcJcznj+UoGn1yH50McsdSGZV2wlXV3jnnftWWRdnVpeaBZKV
X6Ag7k0eDSQzqYgf9QKOSL0VFbsBjIYdq6LDUoM5bQHOAd3NnLu440NRqQWfIhsZnL1ZlSnH88yj
vlT/1lExYQMCmSKtnv0H9c9Oa/X1FYlTitxOXIeTvr1tcUCXm6D5dA5LSEIpDCwbJi34azAO7d4n
E94vNClhDPwK0YOSELGLLfxWAYW80mp8KUwCn68piH6+RUNjDr2Bs3nY8LJ66nUKyognvZhrmtWQ
relsn07z9QFSSCpO1qHsVPwSBPN5vSsL37c15sB0bvH2sgLRDewbNeFaVDZgx4FClwsV2cHsxC8z
kBBorrKal7SOnt1chQjWaMOgiK7pD6RZG2TcrHtzo2YvAoyv50dfdA1t3VjawqM+bheUyOyloSWo
MQ1yQLuIB/1+rDpUsvgKYVAkPkb2WHWRYR1bLTTep/Dby9Is9XSlqjrznW2y7lUPCuJTZSrNypBe
M16bC4gDOnfCjPCOG0cAdgm5LE6bq4Ck9XTPoPZMC8NDarqJNzoV01wq2ocENPcVGoUYQnebn/vA
PjMzYP4odky6v2mUOmVrJh/OChZvTD/ErtNdOpzYIQAHP0snC0LzA8ZMw35Xv/4SvUhYwV8sLOhs
V/ocYdMnyinZg7p2/Nc3W7ATpzjEVzVJLSf4yvQI0sjdUcV5Uw1/XHLcOjU//rCKDw6gAxYpAosf
tLGTvNAbTfKY1+bIkWYKdnf8MXye4l7hcrDj7wfBO0FXkNUroNmsq0nkquLAMkQ6J4GhKbITDuF4
v+uuZw1Yd6jeXmZssCq/Ud4kOPi4nfEVyDW8qgtwLQS93WdqWDSed9bm/MgZE0MzpzPjXqsf4Yqh
D4cK1nvLZs6qrfa+eAMkEz8cW3R/q1ct/4aYkB4Uo0OcoI06Kbdx6YbdSMObtDq/NRFNNbFNrKw3
4+FPQRtlCNxUirqE/Zc1aB/taof9uzQjED3TH3C25yppfuTffX8t+1ie92oqeb7hegfnO4vqBZdp
qlaE4pw7d3clExuQdqLVeLm3FVhTMJS8OBAFgEirD4xAQF90pfDDgcCZftr7RkezAWwx2BTFMdIU
0bnLJu0LB9EDgYCUZLGRPbqOm50gqYp3aiHoW7y0pFnpMi3IzPqCuzJN2oWlwuvKFOF32pejccum
hs+eVyzuIKWWpJPICqHdkBrxLGDmGenEDuB/PpgzJW9bdVdNmPblPYq4iYrYuC9mbacTa+rRZs9k
DYBdtcW1HnRwPcpuTacHXzTve6KzNZIU41YRZjetjbuobHmPC7uZN1s4k4m3ZEPCxb4y2hzfTOBS
qSscTCLlFVWD8ES0wDj9XQ/j7S9kdm+tpG5r38RY3DEhk3cBkH9/6bEmpiJRB4fWU8CE074bq/1Y
RjUQY1a2cpfhx1pN+HSRoHy+P28tp8poYuvPOXb1+lczLPYrgKPpRBUOUxXw4cvFZe0m/H/i+iGZ
YfXw6Z+4BbZ7JnJ3ws7k9y3NXwk4yrjMYlDYaNBzaySrkM2zAHbC8/e8RfgU7Jnh7sNGIer0CjJZ
q738yqbh1xAsi+5c0A4L64aW1bpO6Q5ylTPEBjWRi+7SvSbtp76XNevN4IKH76eXm9GlwjiLt2A9
TrC7LWNv6+xHDffmIhMVGa5uC1Wp+MuOZA6O3Ov/Q2PQgK6NUQ+wdN5FzKV9ygKC1FTUj0ShyDKc
jIm/IPl/XjKVuOvgCcIHvE1Mko1Wjn0TalR3Co4X0xIkBzXTgxEsZ67VqmJPpwIVNvizkdrLvOQv
S/Man30R2nwXUY5IDdzs6qt9SXUUSYM10gVvB2+6w28VA2nS03RPo1Z/cqdXD5eMysLsV52d7PJM
h2t7Ev+k7I2jTfmr5lOsGdwXc9CW/AoAbMIJeCxu2OxZqJRMUaw1XB/0oQi4+Jmg9dOoPInFx2bI
29UOy9+tFJU/IMVSDN6rA5XiRHOivDpDe0viq03ToGZlNIsZnSLbwhU+70vvZox/4Ft7K7XfqBhj
CVZDLDgwC8hPCxwRmbRphP9KHCDTSBUQhaOxGqjj6kSzXhb1rHhSIRNlE7Ue3FWCcLYDOAg7NVox
UNLyd1rRz9nZrEMsl2yJ0RMmJo3Hav/zcWaDZs1YFp+6GVT8ir549FOJXSeowBrD0i34Budd3mIR
DRM+CU7EI1tm14lgU9bZJfEWxtU00tpkpxtLOaK4gCNxWRLtoaUVkmMwYnrx0EgJ73LvK9ap0C16
AFylfPnOM8waxWFkQzE9HNSZWKN+VqHNmBmJ5hn5x6LDSfJiKLhNHwQHERwyawpVS2kCrxqlE1BR
M4LbkdSZD/1WkCQ3iZoUJZF2+pODu0XO+kJcep/IORulle/rYoB9vXtdhoBSN1TWHD2FCgV3UwU/
reef2L48X/DER7LytcdcPxRfnhhUn1x/lRv1BE7pwCvpaneUXuRgaK/DL5OyeQangYVfiEIvuu0R
puFR+YCQU1sqL4aNs/Mfic1SkhyqY9AYUTdIxNRO6Kr7Apn4oogZQaC9QNvmNVbX123Oplrx4nW9
HPI/ajWrvbEE3KdlYeKcW4PH4WDBva/xyvHPEKw7RlRho2Aq0aovF122TdAhMkTRhGaWBckI8UEB
8jIZPQRJvGLd3zQ6QaK/FRACAlRQrl1CIqGHzuMTqGYWDRrySDVpmCgKTGHSCEWGAnYcrLCfATfd
hjlQbpOyLt5l4PT853bOqoHQquxvG50C1Eb66sgs4O0+GKF2jSzc63f+8RTyXyIgU1R31SajhAa3
o0OavMqely8UBoqHuab3ALbo4Fs+PEJYv+YAfGgHWVqNsOXOau/Ytq7MNto3dVuI0lNSAy9sExwY
L4R0AXqW3H9UZ12vZGB6G3jmRcEfNHUGr4ayMSs3s6Zwz+pp+rU8nHcPrOxOcw6dh6lr8Nz3Oa2w
Kmu21rAn+QL1olRqbFZUQOaWy/17vOKOH50LN84gBtseti+2b+R5/nFy/aX+eaCjuHObUbZIi/TW
JUM2gCCAt5uFwFEk5o4hIg1+HFgO7cKraNloR2c2EQnkotHyDOEaG8cMF4s0HyCVnN3dcoZ7Ur6c
TNyEI0jaiOrwLv8cCq2Im+yOuP5fKwxHh1FYd47phWWAtE7lcSyNTIUs3XSmAipTm7zRPPPCkufy
CVF1G3jCAZv0UmC3aqDpyrL2CS7LZgZnBwMtmu3yz06FisXdZ8m7233QGxdQgNtiz/GG6nGBB2M5
IL4fXFSxw9HcZ8LdmNmx88GgEa1lBrwtI28ROS7kTx4orIBtUUHNbs/x9Qhlh3AslmgPaJGW/ixL
oEJwJADbgE3iiQat3ODPtdRWf9vXRG1fXcFS596ikO4mwdty/Bh+C77Q7lLMSuGkITJ1wrjFzcYs
Kblg7U0uNRHsVRzzSPIDAbRyKQg8ABsqibgakqU0CarIWeSZhZz1RzLFpwfc3d7M2aHEtZqaHHa2
js8dglFgyPYCrU41WS6YizY722QLTiv40eW0VnM9n0oVJCxsQiPb5rSKNUgARfPJHMU79nOGrCIO
+BZT92QTMDWidh7rZfm1JUguYbwsR7dw9Xq2NzhGeNpEUGaM0zy6hOThyw1HkHPkhwnEQhs1FyOB
X421wodVeHuzvaDp0abYvM+mNBLn8Be82YBkVeA4Nnqu9pGD1ql/dioqft00q3UGEkcF8soUbTun
nyxah6nAl6YbxPMpzI8ZnT7BCm+pWMCUnUpJmjSKMW1ul5d0EKUY1jua9NkacIhuZDUkg1byu3ka
9lIXizjjhGURoO971GYZcfIcu2IcuBrV6E5udZkKX3lmdo2VcazyvMRx85YIH2o/AfFtRAY8KZpY
o8q1Qdb5xJgkRlCSV4exjA/yXnywJ0EcTv9wqxb+vmNyQR3VXU4clMR+5f8ufNNyusEf3mfBgFhf
d+DrgbsiVIMsfLBLME9S77YFoC0JuiAwmh6U7dXpS35CUuIpTm/OI/oLu4W3AXZyof+/OWY+qYMt
anvsf7Kh+Ho24kjTmA0TdahCXVmYR6HA5HIOSj6d9S0cd/gc5I6OpfA6baBXntavJ6LR7jXP6Fb8
4qkDgOPEHIG4ENvzncjQFFUBLBEind+W17gahTpOVrB8UowWD9T5BceOEgtqbNDy8BfQxfMXWd4J
tjj+Y1ebEdTT05ZYmTDeZ+w1KX/eRFIDAVB7L5YOuBEI1pFXxJfrbRszQ9tLqrCa2+pGdUQ7/b9h
xZGoXyhFaM9ORkQsrGBUMPowHoXQp7jOsAdehqM7y2i/o3pax64d0415oe8iRO1WoTOSQS65yOJU
p+nQjRWIRy5J/IEnHGz/PeSvImNWkCECOUJfUkynpMCZSb7DjdFrWtM5TUWvf/oIQWyFQjIwfZLe
XjdJFe8lqqTt0WVt1fwffyHy46pHqLxPaqhzAQBPeHUgmKds07RXk0/CjD+kNX4uhqnbxLV9prID
D1fvfB+1Bpd+3qJjblkWjxXSyvU/2NGRe+txzj5Gov97sPScfasYj5uTd1y/ojbnQ5dt5fOlQ63r
ddiLIE7gx0+9YuoSrJqn1TZkNP+EySQdY8PwKqAHAWmlc7//Pyj3g+aHOWyUJvGb5Ksds7qQYh/X
VM87WmHiJH9Yfd3lCnWrLZxOMrXguNU5f25kF4oIQntXRAPNjfD/R1dKQdBNWdnOGTBje86PSWTA
vzFyELXvqMAzSPrfDt6Ux5S03ZJ6fWXcu5lVhSC9G6VBEPTfUfZLO6r5bmAQOeFoxtnWZuK9DLc7
tidd0RU1SALtLvMOa42m4PwiN4A2FI2eNencwKiqw2OO53Psn53vHFkLFPkX2v4rUaL1UA0Z6Wcg
0Rsv0rxZN7qQC59UP3JtqWnTdtlg0kJiW5FozbHU9FuQ6ECAN5Ou7GBe2ppy/YBYCWjViYdQXqeY
0PambR+8RK7IieZBkR7541p/qX8mgx3x4sryorioSEbisNxV3ihSwcXnOY/74vIJ+i/8IdxfTuKF
V7bYWtaHa9jcQjaOYl3EqEgIE+TnZuLH1oscj6tw/uwWDy8R0aAOr1oxIxf44ZO8O85pJKwAkrMl
nczqfzsvzzJiI3X2ATezCQBaUj5pojkS3cZpxNDhj3bVosygiVZLWNfWRYTLeKWKAPPqJYa7CLZX
Hj4hxbmbgDdlrcc5i10nN93lpRxaXQONg85Vmt4cTDzO8oR4cr4R84zwVWqmivCN4MZMTbTXWaZx
xCB1m0DYAb72ejetluerFV78HvgpjhzeLXXMYAGy1wIG8lZiEsSmfRs/k4Ue5Pn7+Qcpc58fhNo6
9G3+IJQ6h5kVpLhKJ8YIMpNkzYCAk1Gvxvn2PdKcIyNfYaYoBcwjRNqSus74i2L5RLz14rav36WT
A3PxRGhpBxKcyYCVD7+OO9twQwtQmtoTZKwh1USQhckGWYhi2y4IjndJuAvvFCDI55FJy7x4Q/sY
go08y42WfQmfjU3qnVxQyqi+LsbS6vgthyqCK5l83SKO7lWsJEHmDb6u8CE3JQrlGJvvzWYxd1VM
jrCadNqRLbFiX56xI5Pfzo7AtowunsKGWsI9JwTHtVHQV3mL/LnjD+lUcPjhMTCH5Ze/Vz4KjbX2
k/uitZRocJXyk+7DyqwDUT2SfX4kYtA80+EPJm6TXlnsJcGQ4FanJfJOrDw6XEJLweBYPr8IoF94
6FnZu3ST1nG2Qi0n5FY3TzTEXBOvDVnu+j3KsCukS5Rnx5jlho8snNuW5XeBYpTMvB54dJNXupJt
Aovrj5BzZRs+HqFy/icBv1SkZf63BZa4BVhJB5aeu2qZZz+fiBKiqVemRE2YzZrYB5KBbHEER4sW
nn8FpJqsS2ET2Jyf3YOjzxsYY0cVGZlSfo2GFy5KhPksaG3RprEhnQ8Lzz/qsvh0kfMhyOUhyUtE
EXJ+NnfOm7CEyfx4Ram3ieUuQfxIXb4BKUy5SQ3wO4hWaVhcBl1XJ8HKecyx8253Ye5faXv2VwQR
V1eXDznHC6M4grCvpQqx++l4E8boOp5m4tswojyk/MEj9SR0UjLzfNq8wwi7ylcKF5sr8b2UmhyL
Q95wn9bEn0fydt3hndVt1o8PFjZnfQO7laWmZQ3MKmrceGKDSN1MRwj8OelupD9R9zAtJ9ioyZ3e
hGneFf5RhdqIerIot2e4WOG0rug6/We0Ccg8U+BVHp7PUIZpVPw71l5zEFcSeU+8TC/DzTQna+/3
zcdp8voIXBuEQdW1KZtxq32786MnKYHizKAiDuSbreOOoFZrYliD5jHtcIC/Avug2SkCTaD/o/Oz
vxk2mjNxxDoUGhWCU4HdAgaGrgxpaMTPTYd5v3nUnNeAU1/BYoNL+lr8ll0E2WHoJcjUFV3rZHDz
qZ2hB3d+U5QgQaIOnqeY/HIKsETU9J+P6Uud35p4/bgzU7Rpa+JFYYZGiS+BQ+zR/z8Zy3UPXKP2
qS401pVUWjFD5XX+/n5ibFKChQmsENuvpwiWmQNQQcuwdoUdQukEI76npYp3xiOK2FnXBHndCPTR
/RbEuseHpqshwShVABu3mNCzlp4ablGLeVPAx7H1bcywzxfxeyeL7OR/20hKmN72+usmH0z34/AP
/7Cxe/83T2/nfpgobZYVW2/hzhec7zMmz3NsRglL3U0wT1qwz7VH0l9WsPcv7FmMRqgrKrAk+dKM
fIL6KMEJqZoT5+btCblpqTg52Tww4ecsJAUg8wD+hzYzSMVLs+3k58xgQ19qgzZ4dIat9sCQWxe8
DsijQo/tgQ7M90TMdcEtVF5dksSvxDEzwGqo4fCuDIZoxSImPsaDmtsSx3rUKfx/VMOVjZkI4tbw
rnt7B1nseYZrfIaYKqKAq3oaSNRVKZrZa6V/UF5R28cm24Ob/XoI8mVVQUDpYFvQGfaKWCAGx+VO
6omp1rrD2DBc3Fnt+n/dU4Li0tRm3rCmgD4Sz8b7I6qzx7rCTtxDl9iEpp9pJztgNnrf2X1mmgjo
4umKzIQrQvdlSmtrCeJxsjJibnzZRY7QqWyZYaSWolV1fAXroOCv+lTC18weYxUElvPZgzFi+YpH
noDquHMosj3y5sjUqW3aFucRw1tBqlUcJvYGavekeI23CVBfPWQ8rGgCg+fPpmZ2RxQ7szKPJQxU
vtJXMUd5YYaKxhfsQAoH96dhpKKzWSSl0htf/+I+N08K1oRAdVX6vLcP2vm3gjWiogrmkvFScbty
CB8KbA2cYaWTB+c37neZgPgbFl4cJK0YjwHTZyxKbxoOimB8iJ2tUs838NWz14Xz+fGsY6+DJLC2
Z0nOQVzUFTB3I2lQgPyhjosPmE3KM6PR5/BBemi/g5uITq6z+fIH7D+gLQXshiIeky/YdzpSfAik
FPQFn4QqPpc86TKzX2HelTEm+IWVchvf4CS0VwnHANP5opFciGMSCak2bIhbRcFl2vQVgWhi1QtS
2g0xMC0qfvKXvDsvkvweEPFxIg/8HcHyUiHX+lDGRCh3MBJn8eKHxNHtXdq5FxI1PC4da8G1cobT
7fibRYl5kxcn1sHLEEIFwbEDUueZX/udew4iMJ0E3AZKQcYRmN9AgYOt5zZriTMOLWHpYrHq8b1+
DZCd3pmrg044j55A4y308852rygXGNSfZExgjIaB5w+tZ/jYqJ3WV6WXAjtgGHEDKrX+UYDrUt5s
J4vBDFigCRfEiQuehmWH1NixluLwKg2MCFyATejf8U3+sQt9bmEDKF8giJw3OS3/4RuqcLEz0Wwq
+80hjPNezrlV/d0g9UHPn6Xx+rH/d3MO0ULst+ffBS4pQfXIHKQJ/fBsJeCvIc55pZFUCpUywRNh
TDto1yGpJ2BetuMHTA4gGayEst71e7xz60rWnyD7PoTv12l/sxuXISmZ72DCnx0/WMJfXIuUQaVx
0xEySqllxxsLujJr8bwm7v86jiktAqyjI7AAdrlciFUpwPUthWS+8INolGLD2bwCPdFc4RL0OGdH
KFyMi/IvWDeim3MaBn0LVNid6utRf34ZFg14jgnW6YGQu08LSifvwrXUIwrr4Wyj4579QKnJcG/X
je8B6zEicOUbVi2BFJQGZGiI4uzvPglX5lZwWCe4syZfBkc1lsFkC/I1SKKJG5cVjyFV7dw5n9Ku
tEQ25ZhfJao8kCmDhwsFcgO2W6TN2kBCVIRhulGQKeEz6q/+UsM0WJ4/2D8YsPYm+0VPMwz9+4m0
FephsxAtneknZQk6cyVLW8ftPNGCeRUI67+LLylRnItBgTi+0thfv0E2B54xDI/7mGcrj3dq49G3
QsyS7zngpYsfS5uXvQkvUasarpe7aWHk5F/12x338n080USNQTrSxYBceFVCi7ske0BY1ou7ln93
vXkihPac/JkThqZxJTmI+tJ0lY6WYUy6Gqfcy80Sfu7Z/YHt+nK+Ehf80UYCjkw65WZsr/xfxbfY
1bB5/5zmGMmt1HSfrQlGmqUhc9WQgcZyZkvawz1iiWAX61bsNv7kdbW6tqtBsbk3vx7Sacln6z2o
FlAo2i6FA3Mn/4yupLG+Jzc67Yd2eV5Q9Gz3+Ke5G9hAWyFcnDnujPH/VDvuAst3BFx/Y4tv8QgY
UzRAWLSZkQ05j8o/RYwCyXVsjK29YP/6wSOq5b+04NkYcBQmT4KeLWW4jEEjlKTt5l3ZVerRsPe4
dGkBfTEjDfJEWxO8c5mMKfDQMdh0hsSHRerImA9fcznj4CSvsgewpjicDyZd1nETxFqwiFeEseL9
eoHnkdP5EaPoz1DxXCWV5mXHT3VD2sL6XS777bZEdoXnKh5wB9Z8I64exUK10LHADwv5Bp52fu6V
BFZ9oichJjNhfatMMr64qQxjjmWqMUSbfe34gZMbUfhK1/J0e+XLCkGRjyaguujzJAEbuAX/ZPha
6FLhGnSuIb/2ReUxLRMrtxS79rCnV/uSHVKmgzfq4RS/o0CTrMXwbqRMHdLQqcgbdK2qk6Wb1Nlg
s08gPyWowT8X7ODADHiKQri8pHZpljUyU7wldiNTW4oA52h/UShxC7Z9Kt4Ewa5jnkesL8mOles+
ZJtG7CEUkffSsVu8XDZ9/VWbbaCEKQBTn7n6et9lqR+HzcSoJHqVUQTJekg98J9pp1K5iHCIkYqj
Vs6eMiuHaruakFAU8RSixxYQbnKobIFrEt6nOfAO2r2OdzOgyDUS2pWcFk/iH5pASsrdwE9WyHes
d3GJFw5m69ZEdF8uWp4pZMjwzduf/ByNLNW2bhGOhArBO4H2Tpi8Z9d2RHL5wZDS0sy1osZlnI/K
A0qEc1V9pXUZ1G+8nb+TYMViOeaNpWTHHZm44hrqnDyLgwfuKjZHeqYJqHBgbEEFRZjFnHzantLq
YPCsSFJ65YcdU39QXFBFkV7KSyfUI/fatRuwAQLaizv8AxsQ436+v5Xykjtdb9kymA0Zq9ZgZKeH
DunMU1HwSNAxhVovcdMKJy6bEqSwrg5lByKZOYDgjTILCGs3qXyZeT9g8jl50gKvTMicldlY2SjW
/JbPZaI5gDG2mH5vndQWKUCoE2Xt05x05ypi2776MosqfYvVkXiwBc1PukEz0MOIjEIyqe2STlJf
1gQF3Z6SlBDCpTxxLpMLrc8gk3n4LyVrVQ/fFlG8QUBv6QHi3Y7k9FQCLvwLdNYQXFZNEs0VVcGm
XW1TIYd4z9QqVs9zEw+lAI0vKYOB442h4J7pgv99UqFfM1oweOGxTQurbDE0M4o/7eHvMHt/5Zhj
9BKdTjYthuDj1OPfYxf8JndvijSDqQ0MOHKGhHjwaDY9G1gzEBw5afgFOlEU+sqK4WdHE+17pS6F
LkoZwVUQGJGW3plNtT4UO4B7tO/lN7gjbOiwDT2lYrAq+fz1IN0Wqls6N/TQC5eWikNAI5j05QFh
sJ8bZzjk8XcUG7z37W9hzP3qmZDXdrLoV+mlneu4r+z0SLvzOivBfjdJXk0fzV3ZGQMy4KnNRJsK
9OvNCruzlRGTmB/umnRa4qjRxMqg4xd/EkTFtY9xQ6BjP/msSDsorbOLmkj0k7zqFXtoLUp1y+DG
ICTRGEpZ/pGbRMUTg3oDvkozONVQgSJXwKAfRbSP5Th0RYXlcZ0L/qc/BrFcvOxQHBgTfQsQDpWb
tRWuc3chTXPMtGoqQz7vqsqPsNqMB9AM8APKryGKYRnJeuOsYrZWjQaZx2mDEwZ8+4JIEaOpHT3T
Hh/9fRZcpTuwSM1pbeLTWTKPh/yzznM2sgRQz+aXTC7B3fK4LusrlRVI3ZUmeLohykpwrUM0rbm6
6xPcF8y6YZVAa1Kz/YSlsVVNN6LoGB13I8P+X3DPoTpsvgx6r2CV2SzkeGpgKM4su0wBLTvoJCBA
gWFqBmsYlzthWt+KwIl6jIMY9X7LdOZbsiZGAnoN6UUKb8LpKwM3IqJDS7iQ39xZwjy6oRX+eIKi
tfT8LTdVVce4iEyAWvKKedyEsFUCt1TiDRp/mdF6bV3aXKgNTBKoqfce5I+4EZgY/UOXsxb+TRI0
MbM+JWk3LKazZWlCq/MAfRZNzLznNhozDCe20O+JCNbRUfsHQWyWnAQmawM2GBouCJlSjFjwCNgg
uEbMoN1WXVtrTY893uKOzMMWd/p7JtNjDF6VQ9cRX0dc4RUfFkSkOmndguErODvBW0pMM+Jr9I2j
+L++xUJ+JuKOduwrzNrdAF0PBHyelDFlFPSpdQSp9Oczo/KV9owYasobyJ/e9XHEQBLrDt7kWyuj
te/nVNKKdROLaxnrUfoqNpJElwXqf2eW8g3uiZjUxwAeDny8X6IX61cipM2m6VlJebhQJM97nara
/aPu+Ow2rxCvXcZH3qUiRPuf8SKm16AuIIOamUCtIHtj3TQBBIOvvoyXdDC51rwfjUA3uZiLDqVQ
d1uKjpSNKOo4H6aVA41YL1kyQCoRChhxfyqvXobv7WjqLvDqJm5GP8vo/FnwiWCNeZcb8Ej9ZpQu
CGCM5XUcCh3cb4vqB15lWy4vJUBGIjXiq9yQPppfEsrXOUcSMZN7j5PHA0hbeTMlxibM74q6q+ec
muCQyR6gTLRFuLrMqpI7fhwTe0Xgo7Ab+pbLvlA8nlfw687kcvutP2jCnPd5WUOqZ8FcJla8rLzx
lnZsKYxqILbv59JyPZP9rGwz9yf7NiZFOMlXXIna7zyjel/eHWlkXhKkL7kZl7puFCiVQ58Wyb9I
IjuK7vX4ux4bJSu+xECf4187wcnj57jPFO36AYeoscPIFr9Vd1DJm/M73BOnYSpOT3rgzt9lCTav
4JX+uIOVxKagUYUVlaLYDNFcQUPKQlKDJn9alx3OJ/epfplWIXjclAr2Ixd+D0zU4nI+J4tDgm1Q
dtq0RXrYe/KYv6uxdVUUSr9FNprKhaLtX34DDMbhfAZbEmrHyGJ7BXUf0zMT5DM8SCUm6Hp6yk/o
lz7CgfPZFiB+cKzbSntAxTPVb8WmqtfGsV5BYYIHdslIkRRmWHlGOcuJ8o48ZLjJzW+HwuHDHlRR
IwDzae5T1ycV3yEubzcrDoBxMRO62ieCSgY0Sg7M9T8+W1StMWEMG3cKsmrPBU+SNjNYoFUSLk6C
0fBOZ5gJcI7s+ba8tgnktce/hYVHmH1iDtCMFcrSa+GbJFcPf5xIxxiVMdKf298AVgU5zDg7Igf8
JwSFOZiSzNX90sMqXjnd3lypgqINNr5BNmQ4IjqrgERF3CbaL329nNV6+Ajxb+NbxYzkOCHXkmr8
298nUxvVUjkVbo0j5jLrt3r8Jvq6dDjtwjENauxmByyITcWOuJBcnn8hJrqgvdrmjZMUsTfgKaVr
hbXQhR0aLkwT3sdd9wS+fCDPYEKYXVfZWeIMd2YhUIIkSIZHWAGEPa/cj4cmm/qj4aQmCJkptYBq
4IfYoe+yeypJZ8AOyi75cH8SKiyQ8TuPXHz0RFGeS5IrTs4XuAT9SbPSTMWv1BEfRqTT7GcpBryg
bgN8ub4w/ITS4GEk5ge3IHn0a8XHnRUs6w3Ko8dE5LUCS/4U36KNIqwIJvgRgSEP6odQhYBaCZ3R
DzvnLdKw934H5KxINW+5FO5TGhH0X4yuxVwmn44/cmYjwbdCM79mYKD3ZBLn02s39SzMYLPIFpLz
dFGhaN04EMI1KgVBOyFfkBKpgjDKv2tdPIICSsfWH65q3bt9m4vEGv4V1UUG1YCPrmylRU5IWX+E
ZeTfS5QhWW4oFsAzIPghnoht6I9rWq3a2qsYEoeKesz916+azVfUBaV+xpMyMnAHr3q6OVwEyLNG
r+7EQU5DTRQgUNDAGIpye1p4gzXV+VVqz5h+MUhh2kh+XbNuLsZZXTn9ydpTRPHvyAVncHF+kqIC
ZNqdSO7YEgGLrNJxsE5S4IktkkdB74or+/xpcLuXsRqjChQtmY5v04GdRZcr5iFvJOr+prdvakOS
EyGY3/nkXBhYGHV7ea/qUizTJFknQroJ8M1QEZkLMmYheYVhutlG5ATaoVxoVpEFLRY5RBz4P6c4
8C0Rp7fCJIHmrwh3Xv8oeviNg2GePVf7wB+ZYVIUa4Bg9ed4EsPsg4vdss/yPXwvVSqGwJtljZrv
NMCLjpi7Jcm+2nWeLmwKd6kShB2CRqUnKnj018X4u1I1sE+TJxqoEtpdVReF0tfu3z2bt4L7nuuu
hNweUjePhPpZL7T1Q8VRHgHzxHokzzyXlLPBWuMQB7n/uHIUOTs8EoOg2L5QpLRgMlcJwgaVueaG
qYgSPsq2pguy2K+958RKYySNs6uh0JeMGsHipXZqs6aGeg7sjIIDwjjoyfH2iz37AXwY+XisTxLh
LmhpzFTmNboNGsPYGSoSvfpXMW+EN0tQQVaqfW1InfJppyiS1GdUZd22/JiLjJAzss56oe/luprL
OT9pMOUmLbH04mJGHXAUAFDRN0zjv8nP+NhYQP9ETQbmhqjg/zEw9I1HgeUOYJLnbFVSUQI7CC65
sBNGjNe9Ufe7Lc3IMuNXEWUWbdiDHCqYz+dbPGUb8YNar1lZS/Y146QDsm+0wdnQeoaxAQmB1lnf
VuowyJB+xq2b2aHiGcByP13MBEQUSbtCvy7fpLjVfPqi7x3kT+zy8d9rmqAUdBc32+r753XUfOA5
+tT/FbMGSPIhcvcxYeR41TV94G74rhfhbBmmjnfCP+CiRmku/Pby/0E01mvVNQXx2qdanPnysSOt
93oj5zamvoS3oHqBOalvl/GSAIHJ2YR5xm3CHYSvyBoJQnpnVgBA3SBYIZ3Hiaacb4SqbNpbtUKm
DOVgDy7nvBetWqtXJ4qKhq5uzPARG7qdj3MEmVCL7KRiIyWnSOvZX5yUQg/QvS4V9T74q5MEZ8Px
G+EsRnJUge6+2imMjBUvOdmH/9jIlJOlttkqyEby2V1dfoZqn6ieXzpLRYHOOgaCDKisEGOJwUzP
z4BByoZrfBjF6qSuoCCu3Dl+u2DdAwJOyG0nyjk0tl5MR/JOtduwK5meaUWtaMi2LAIxQl2Qo+kM
C/Iir3WZqjS3hd4TAqKDhoTMdso56HUnSmXNI6IvEff9Kp/hMtYi6KXcjawJi02feWCMfIJTTNU3
M6ihDCbxmpX9yRkFplJVHwYTuQJnmIWkNrvSxA0updYARubOIIY8q2MMFlumdpV+IHtxuDdrMRUi
JqP83Zr7uHI+k7+jfy89MaFQJTlp5Bt7i3tW9spmImnUQv3w2ROgIlthAabavbzjlDg0qPO1BIzD
aIWsQdenBDa/xW8uGXb+ZW8tHdYcQ5eF5MHpBQtIgIxRbpMbN4B8XxKx1XtC1GQGv90n9rbGgQGx
SSol3yVxWoITh6r2x78iVnu9dZgYmtHqbCdJXdxhK6PqdtNzsITuzV8Qk2F1xqHEGwZEbs1NVr87
q/ChFDHEpqLIhry3s5xBTbaKMXrhxDQ4xZ6GGEyRAAYebjB1k9NcxYC4jbUphzfifOfMt9Rn4eqG
Mz7MDAU7FmOo7/ykUcawypwDUfMcKIZCLBfP1RgImafN0dDqnFvHIyg8DFFF2klpcw4BZlcm31T7
6KTsgu8TbtZIOldswZlodMrWojFrh4t9+AelBslGxsIoDnOycvfKPJErhWRPMakJVR6VtH4U0/ca
Pv2FDvjCjg+/61z11yjIHcwpi9PI94XDQPxmV9lrng6hsvNlORLD9Qu6Gmd/MKfmWr4ksfsDAKkw
/oFsHz1iyqPXj9KyfF6LiMvWB5v4GY7L2QjtsbqPCVJbKFI5oBZMZSyJDhSnwKqc7rH1H8b4nf0o
hFxOz5bNRJ6eknRAXHOHcduPb1jkqUoRSYaHzeeq+pPhtjDq3qLO9wBKILb1xXzrFCpSCOAhZTNn
P39YGKIeveGllAO7rVJbOcCUB8bNZ9dLJtjATVi/n2iMh9xPh2edXqZQQrVQIdWlxudlpqFR2Igs
r9gRBv+dBP7UOWuQnRYVRDIWGgh7ut2pyhssadhZ9MkAYrgPRGTGt1r6z3x9ui2H2uO+fTpIUuRW
nKp4ETWZerSHG1h0nWFx1eCj68OlagpcwmJX1+2aMPz31cW7rh+BigPoTQqiTYy94q0mNVdxIFCj
uIx3j0E4VBt5PlhFMu+gxDQhBswuzrsQzLl6WQzbCN8oQQO/nZQ2Ml6lJXuiwPvMdZLeEZUs9kpQ
AuLCPjUjZDqo3K0VR622GhIiHXPaX5kU41rUt+pesXNk59jqhsvkMl03ZM4m8AsyYm9vJInc+6pf
XO9ktPvnQwAME797ZDNHjagUJ7NixjtASBstuiI0haLM5jcY3kzaGhy0UX7WEAV5KyzE09hEupf6
Q6AhXe8OrV3MwaVdc8Zg3MmCWAuQR75iWRl7E2vUqa9a1bKHZvAtDiJVQ81x2ugpVRWlI5hBv3TF
GkNdJ8L45DFGhMdSbGt9GXOantGkD3D8kYYFzY/+pdR8XT44W2ADPKjxV9l52Gtb5+Je1491c4Ox
OJ6U3GFAl5Z03CLtxnXZ9uXftn8YT+FQ+8LquTHfJrGKilGnpJNwTnc403edlH8jZ9by2W5A/ElB
rr3ffGNUQVidqwX9bSdUYAI2ZjdE9WhCu8OEsnqT0UDvMLHO4xNrhgle5HCl4iDK7yobGxIAlpXg
LSjrU2PAZqO/PKIaj9cT6kOK5dLeCUS/I2ToeKE2I/WLkg0fZjhyc6OgZPMS19fD+KtfEgFaoY2R
djccbNQp7yTZ8bIFWmfkBLlimgjU19Qvh0psnmfFinb65VIEkb7RDEyWvd0t22BA07ipfh4sIkmM
Lqtk1JSGdQVCiTdCQVEY4ftOPYXSRaMMs1VU6zc7dWsfDSCxCirKxO8PkACLtabb2vl0gk+Ur5aA
79VwZzc82tJPOzZrG1rez617d8xfEuL0wGjglKbEm1ypV3wh5XctSqwdzKVA1jwc+20UUwcr8PBY
HLNIfNCjFZEC7ya+5UYlDn835nNcI4Q4AekLCiOyeFPGlRPfY7rKus6XmFWlPOkQChU9Bmv40xGr
EVzxc6sG7InpUHQP2BZWSae/QWDTgnPkfaCTUnalrdDnxH5Vh+nygVfAjN6lv39uen0nrOO9wbRl
LETRuecdHOiT5XNlU15YwBf2m7HhTic3RN64nKCE+up8uPEfTZtCeM5xLW0S0Xd3cSYzwmQZo5B2
MEXobxhLxCM0obLAQEe6dHW6rtpGm9GYdUbjsrwAlKkLIIOXJDsvzVqUb1ikQuAAekYH8ie9bFbh
EXloxYr7JxxW8p5AIU4c1uxfrpFtXwqiQMMoU4lWVZYmkmhPOkWGmMgho6/INf47UFgkeApFY3Yd
xSKedYuxCwc1ikX7BFhH5tZTp+Gn7y+rKFrremzk/+V9RldtuMB0VFFQ8z+3LXEAi1y8LIGMevXn
YGljBS2RZl0W3FUd5PvcinyXyukoXYWy9BFpTNfvBKVyEm1tmVeR/RI7YG8KObSa629XwELBvIaf
uayOj9PC0yawMmsPOr6fipL9vcPD4ejknaC2xTgTH3qFXo2gELzDbABWrKNUhGv3bwfZNnYDljw1
a3vhqgnYGpqd9OXGN/q9vvDqb4f0d5OCz1gV8Yn5cgqe9lK1VNhZT0MUutDiJ+7UMJIdjeg8yOPO
R0XYFr/sCIDEza6q+1UzpQ75TQe3cwPBs7oFcGXPqdtax0XrSc6yerNdqDoylKjRqsUarXLcUa1M
n0oBr88roB7wTS8t6DvDJOkKI2I4cnRIn5c3imSzBHIUDQSgXkbSniV1KtZbzztm5SX2r3wN+BmM
NRVpThAgSIm4UqiG6khEPBcNN/y8e3w+Q0aGxyIE98e+7uQD5oS2y8oMkhsYoTh6Cl1ScB+Qofic
QT5TFCvz5rSg6OesS1oQWRYdX3Wn9KaIWfRarvGRJB2JHs3bwaoWmjsmc/Wj/TU4My/ukabsWlhT
+vN4a4tUWHKT+ErKrSOtixFGk3Y7aS2Qo1HVYmxDxnbfp/XYh1Cup0JXsdQxsOV3ZniEW/dOtkBY
jMZk4WDE4stwKeKX6KM+PAldB5UE0/2inERr73tk1nLoWWM2CUUXMlhrS/n/huZT/Drk8177vp0x
s8q85Q8TrYTsLOrZgbMvdsCeJMsVbxP0a67T41snjtsYJ3BW7hIxqO+Ej9e+YVYp2yQQu6MmpWJq
iT5gmPQmFbEa3ReM/e2W253EmmIBjNXto/+j7fcOvwTo83vDwi77GKDvxjtnno2n9M/gf0co41sk
sSFYhBgzoAP/iXyDOqQhvVrwVgtFZGMfkJwbZvKhVQxQtPb+7TWIqPfM8UAf3KRcHqrWNfko8T1q
aRewW1EUZVZ5r2yB/i5IJSwy1ELYlihhtwqHoJfIUB7FlRNTpqO8Qa/r6cRkl6y3d01RWV1MsYpn
YL8Uz7cFQgGf9Sr+HziBydDPSgsv3qMyHHeU6+jTc9FHHdyF+l14y54MIIVF8oIkJyvJuX92a58J
LJpgb8yzc93q848QLMMP4Ls56OJHuYL4/rwYu//21MZ/0xOf3FVB3pnOsvTGzp4MLSq7XKet75Mm
yjiv41zaxExijHGNVuZgqMWoaz8+TkHEEhxBdAQXUWTrF6n8bV+qAyZug5lkVecWVoLurS7t+ibw
ceOlXC6n0A9UBCzzfsDruk5XCk44+rHdojdOK+FdA8jfeWTywSWLdGVFgV+bjF08PGt/THXo1wDO
TIOMOugYq+tXO7Vd4Bcpo1q+vm3ODvO+7cdmur3Ye+3Qb050DnPJREj0jYkiTOn0LDOIBeAanIZS
6C7nLvQ8COngKYJekMv3dUTg0+j6avh0VwqE3K0K3vNO8mGA+SnYJe0aiVCF+q4RMcfdlOfUhOIN
+r5xrXFG8XYE1EuJiHp61GDlXJrjMaaSCfaQoZf9Vjyc0srHLiuEsyxkgsf1Uh8+oqJm4qQ8NLSs
ATPuT+fxAErSdweSyWdae289tFY2IQi7I7SA1drWQXSrViKX54qT7h64au3Qg5xrvhRY6EQVdxfn
tYhHG0dfSYYc6eMbRRB9lKwp5JCH69Wh7vrWSGarZ5UHPHmymxpgP6lu8s5iYa0RXDE6g3s0CyPR
gyBBwWvCZekcF4QX7hUDNGHsr7KDGCgTMNfRv7Q9bMm57WZS8Fu4m06R2GJi7p29gbAxVQn4jZyv
rKokZxkeZUI6C6Zajc46qs0slQcj8yXWEqsn0AVW0g2LOAaZ64W0fnAX6rAFOnXYDg6ynw1yyDks
0BaLmVvvEkx/8aUizjf9mquM+Fl6XJ0nYgfHbVx9oDj5fH5PID2j7ExXSxDQC/c5Plrrf7ZObrh3
lXGiklfhDjs+VVGWCMD9uLSQ8aXoMcfhZBM+XjotGmP3Lbl1t2ptp6wosyy1rutC7fIelQ+ZJdGS
ZL53j6xf0lRfvJMdgGiJAQo9dak9yd9ZuCR/94HyiZMFrAI7Y6Lr8rZhZwFWz7roQkaCkOl9gOps
H40nPq+5B41qu1AnFGPJKKkhjsR6Ee9Wn2jSV9CJEVBqNiafKa/AnxUMuS+A+t32wNwhVS/8Tm9x
VdQRO9V6WE/FJF7rzalbxjvmzJ5YcdT2jF/uILNEFrFOGlCnWSDHOkrIU22EVKxHX34hAPHRTYKR
j0QzwtRhCiSXaNbfjJW8bu3JY9N8eu1adS8QwfMChvEIY8BFqrQOFIg3mu3sIYUFJQpQntXyQRTF
Mqy4kEVKF/QdJLcKHWK/VuvYm/KQ434hS9DgpeY/gaBlLTFbkWXPhAsGLXcYxMV/utgi3LGHrer1
/iilVbJtTsLCaDi7s45osvpHlDhOhAq9VvMBziJu6d5IBSAldiMTY5cZL6ksiovMWlz9nsJVnEf4
tFVUvuLo/MdDzc22Q8ysWQ9sB0O+Hvu3QbQQSNYG8SzY/kaO5J45GZAwak2kwJtBUEGwlS+cuE8G
h3iBj82Ye+XHy+/CR0E0SIQiQ8TNxpD1KbK8bgXYTcvb3sVF0C6wq98sQCeN4w2s/e2SVQJAJ4yg
QSMSBHo7xAyZutUL4yjGqSMNIqUpu/0bAg97H1GAbA6OInbpSUbWeN+G1suWjhWMhXUPzNZHnMt7
VhGCHqAgEYG6XIn8RC0TtkCt40nPMxo7dsOUErQDPvs/SgKEio6mupDtH7Tak4eDW29k3HuZN7O/
iudUtQYk3OqqDdi0ihE5tLZNm1uEZMNvxSTw+Hj6tDgTwvVPt+LOQotX+nx7Gv8L8g93/iTuvSki
adp3S78DImudcCPX6HB8IkyxoqHB2e9PMa6+EQr3Fgy2QlVcVC8ixXEPwWSfTd0lRlYGGL3dNRfH
1sW1KowcSxsEj9rCJ4fSz78T+g6mZRqm0UMUkey2tv1w7vyN5BuuKXdtfSmgqzjAuS0bRr9ZD4KM
HBl5JLvO+ETMF3f7HWuKEh/rbH+uZM+xSh9206WpExngO7PQKwEDsXNhbJydZtC0qvw361nvU01i
wFpqL3E4+wvlUEToE//maO4LWnv5v4OFZg6pgrUo8cNGZZcoohTO0jocbuH9rGCqeKexqgEvEPDw
BKMVD+aAzcdr2h3USAabI+mIFoz3N5mzEPP7V/XUmE+fahSKDo9j8lYVRovMJq4o7aHQg3atxJoP
VnFDiZt16rWzyN/1lErmj4jvXpYtTJpnieDpzshVAn9s172BSdJxadTYjfmu5QVqx8aGKRiHHJ+y
RYVxtUFYeXa3nUydYamhNMJl81fg4n674bsO/I2O0I7XtB/eT39+mAHOT3RCs+0P68kwiudTwMre
u7qTZvbQsBH0ol/CShumKn1aURiRHq88524vEpMOExyT8D7er/qMk2sgMRd0eq0rJ+kAKyZDJJnG
7NSoU9tfNS51e7Yn8AtWFiKuum5IiJZVmUQFgWw3em5910YjEF9e0ZkNLXbCEEDNo3c3GipdLUG2
Wf8S8HCEeGE0K9BGOTY3dqikM5G9bz4iW7YfKUtMR0r+jwURqiaMz1HxBaqhxVy4unpNXIii6TI0
CjI7bEEqHuR6FXhUtrdatVbWWiaWzY2sQdFF/giBtH/WMf8CYp3gYMjaict4JjXUXylTXQeVyDEk
YcAtMqBbRBhbbZRd83hCaYY/aX090RE4AMO459DxLGXBFPnZRsRHsLVknLYb6GPE8xHLGWIba7ZS
VuF1j07e4v6juq5SpF40CW6+8tmkCajS2KNOAghFNKr4miQrR/zDepVTLWb4IE/Xd0YwaeFZqaX1
RayW0Mf3Q5XY/BIGD2Tt3ww3AjqD2EGaAoXyUiM3tzaV5Q3n9wHYFgH3yJnooOyQYGzqsjYlUYGF
3PkeA3ZENLXfaMYqnNDU9rGTQFh/dTwyXz/zWyEOhQWZpRHK4kxrx49Ytc7RamSlD/KiZBbUmK2B
FJR2lia4JcdUdeHsFcShDzzpPxmU1sDmYv6UCuCC54OtbxmRPqkkG2P9c04p9vXPw/Q19b+BqF0M
gi7fs+qV/q1ZhX7N7EyVVzQ2E74M4Ifo12QCNkOPjTmNDS/ld8Bb8yiQctd378N4EhS0VxnER+GN
HTn3gopMZX/ru0le50TkJEKToaIgtsF/WiN5tgcf/PruiKw7DcqU+gSgW5zg/TH5GcQ/AT0LhLbm
/nSGWf+a8t6kpHa/xzAyDItYb+ILzzNa1xUctaJzCq++SAoDHwLVyrRabUUZmaaIUT3puJ9SV/e6
JXrAGhdjexkCQsMkE6mVAHe5M+oUgquzABxWFaXn2/k9c20nFCeFJ2LOmuHvMQAWfZ0DWH9F+gEA
gZoBoLyWXIRog9AQyo0zzu2MrQkwUGQkYN9u3VyMvfjLP//OfJ+JYX3SVZrqQtRUrqhq7jmn4Prp
os/MjfbpS45S7Va3Z5qvDMtCMWGFUiofDgTMehHpMKKo8Vr1p2P4eJQ8bSjJOeRnmYuTqrUV82Ur
r0Mj5j4pvq7VtLIWFYg49H2FbFdZj+sFsfaBEwVMtq+xz3FAC6eKV6PNwfiNmv25T9uXjwKXX1pt
Vh+5Aj8BKLrX85HhgZHNQUEQ0ZTBuQErP1WbS2DBQANiMzny15oMIiJzCfV/NFyrqQ871hEb78Jt
iDQN+qfCPCkSAWy/g2ElE/JwJ4O0KTekIyTpbpPR34vbNZg9y2X/v/degpnJKHTy7KHDGT2rZT1j
YCDfaX78t2GzbAuvYFbZ2sYMlmX0Ui0WO2CPDVNoV6rI7OQgK75YSh4QZjvu17YT+EDSngv0D2wS
PXx+7YK77oZe++DGbxJOw9rwuHNXwmw2redFeudcLF+oYYvOLK/ouq75wTCXwF6y9ee/r6rj4REl
WcXZc0H2x75YyxGE3UVEmNqGTD6I9Awd+eiiXYdAW5OicNtIBDEhWOvBQAWgQ4WsQPqWrX6zY98D
0E2Usz9ZGI3jF6AoKV/HOr0evhAYehuS9jFOEqkPikOEbsry+Pdw4EL+moMWR6ZFH4t8xsrAaDND
0CYT+uCewq/+tErGEO50mC4EW+aKOWNYG7BHSzJT/VppKnfmNo+b3bmENjOfu8V3jcKaPVJ5ZFSr
p2RPvUUdxyFPX/yz7RAJ53/u6ruyShvqRJO8W3n+ZXmPL944TyVfYXIonrEsqsAZskNMmMRdBmNF
zJsLuWCKUQiUBk2rkzb+3B7fm4TtPpAfsVJZC0RggzQJ11NDyfBM6JZW+k2O+01XuQv3tfwugSGb
qi9PUBq4zU2jELDAp2wO8kpa2o1+vVyXArhWHygAH4XsG9DkVzRJhUh6BW2zCJJKFPBdUu9QJHzQ
Rmfxw52NBhbNG3f+PcCDqyxpt1Zc/kc7ORvB1+cuyJbGaiGmt84TMpb6cYrWuAzXFRO7HcHqtpmg
YdXUIlLPkR1oCJYlGmTYXpT32UpbkI3vtvx+WerHzxaaa6N7TUfmZnCZBNmXHGtVQxwe3I4nZHa+
sD6laW3CjXCOlbEZeN4K6GAcLsHkjRu+0eDoJMR8z9XW+JWfEi6GlP9w0d2Rwe87r8XcNlnF3d71
LmJg7Uj+mXBJknB/ekUJ6Z05c1/xcG4F6Af6tDN3mzNHxMjHL8BWH67IhIQmWZECgcQvtp+tNb9r
RoyLGHCKtxuzurMWTEpG6yK8aZvY4Z+ZmMgatBPkZFLW/kFeCRQdslgDUV+doRaAd+cMS0oCczRa
uScdyt2nH91WL9YhvhLDMtNwEHbWGARljH6fLHqoORlbDEOVsOku/pEsOuep4m1hFJ8MHju4V+25
OwtEtXUxpBYAcbb++jrDWajYcXz3vLWA3egRc+bXrAtQ9D833k1+z5VEUvhddPwzQOSE8lXML6bg
JwDP+LHIYlXlzNn706dmCrrQEDlUKABgztPYehIdsbt0fwC8QEnvdK612z6jcXiOAqB7H9Jca6Oc
PPoNbQgJAlY8d2W7tYZW+4BNnmXUxCB4M70XL9HTKUiWMNtly/O26hShoiKrLpLymf0hOY7giHjV
hB1eS3MAJm88YziYVY50Ofw1MjnZtyJoixvUk8yhjr2xwNPXdyboUpHLwKbuciId4sK0jQCsWluE
HuhkXLb603dpvXFGZOtUUqL0dC+pOcjgxU6uCSItpIUpZ8rvny8028NqbMXKs+moQ8NLWZzlZKg6
J4dSHLSKIMOF91N/+/l98lkoeYG/LAr6VxdRzAy2SYzgBKr8rp+UczRzgVxHRdZvlP7Cze0/HMXV
VAzpMOexiLnJyZx7VQA2gqjzjE6OypewlEO1ArX+WsjEjFn8AspEZfKvrlZZSiRuxq5e20hFHjwc
e0qfsRY832vLysiuIkwSMgDvC4aL+RBl1nD2Zttj44ajNm9xmfwnKmHtOB9SoSBg68S2QJR8edY2
NnZuJApbOvDdfPviyGnE4cl59ha51PDOZutZe1rfxxHBLE5KxGtJZTSQWwZecKCZDk3GJ0Ln8twx
bS351ScO8t8m6zjIJdKsDkNpWo6BTfHtuPtBMbEQ3WQE4q/Ni0jie34Bc1MEFgjlKmcUnKUpvlzH
Cioxhg5HJdgA5HyJc8XTiCPtX4dcrtb1nq7ViyD5Rj4m1tBsKEB5zpN0u337BY1KONmzG4eDjQ/l
QO1BQxud7dgbLDC6F6dl22phXgYmhOtSituGld6PESf0Fs+dXI/d99SYa1GyzFSWeBYyx5zXDUt2
IJRtn0bfrRthCsK2O+L65RFaa3M8HpyvB0Gpn+Z28S7pFYygC26W1CEiriNsQrsCTUOC1eF+mWNv
VA9hYsdIY1WkqEgS3F/KrDsJVOOux1CYKN0ZW+aZn69ME27eQMQ+3dPhC5BM7O6NgPk+DlzJqI6r
ycSD8MgH2tXtma0Ao4PW4NCVrjXjCaVB0gf9Kg0kq3uxLg+OjXOizGLfWwCioJIf83JvdzM//D5N
kP2eNvAYXeJwwv1LeANW0NOXJgpJv2TLReRVTLfHOleLV/yOP22PwrUwirJI3RFezxpsp3OpPDny
UHvLDzEMhmFlCumgKXvlCcobS26lLPi8+BMJavNL/WWsKNlW0bBtR9n3DD3C1y7eTO4kKGEPK7Lj
Xr83irz8ItAzhASrnz8Gzrtuw6Ex9ZoCdbfV1iX6LF0FztPUk9HGSbx/QQylhaFoNCtZ2Oh12PvF
VCh/eL77igzn/q8+I7lspjoUWdPHtYkAKEv3ZW++BL9X3/n801c8HsFo1VZqTqeLisEEe5qKOiSz
UobXSMl0xt+6BQv1YfSwjmC96CtaFDBi6cYWzPPyYtKPELKoy9i3V5JBq7l4s6HWgM0lo5xL+4sq
78u5y/wAryrEz0IUnnxRPXcoy8bhhM4ARESlesMrLdm0gLtW64GgiL8utrTfYMuCGfifduvXNBCX
RCsJ3Bh9ekJuWWAbYpxl2nc50o+ceE/QmEifWncZTHwMqGUxD6o7noxGz0XGLujGCOM8fCkqrnRu
66UPMpUH7Zjg8FBMSucYSzcrTR+ueZOHP2OFvL8iexOOl80Q1kd2ea6SYE2yGnK5Yh1OVqeWbyIp
XEVCZzH+SKLHXALaB9ljvVsWDOJqOxf46P+64BeJECWJZE6Js36qnff62yZJPghdZY55EIVkGyui
ZobwzRhYAfHJZqvq3MWbhBX/ojfD6wdeDaTqPePvpd3sq8uhXBLng26KDOJLuV1wAPr8CKGcrk+Z
Ak21OHmkt96UyLYeYGTq+ZdGTiBs1u3se01n9vPlbzatkY6w1CBC6H4srRXClisUFj0Nk71ZrKZW
mX9OBQmwxLHzlbiZiU+Nm8oHBC/E72lt7rWltdVrNTbe5G9yEGnVYK+Fg+G/WF0P1GObqoJ0ay+Q
LuvUNOpeKsqtdnLDzxwV2GPwnqSBuXVQXCwFDITXb7w85X4/3eQCamGqTNN9zW/DRre2384RjmbA
+m3O09jpNYeVl58hoJvec+ksLEjDphhZDtvWSvaOgfIjM4UWDunrl9ugLnpQBVb+17ZjSfpfI4iN
pIDRaz4sl2e+tv1tfATK5aYwthuV4+uNLlNcvJQtzpljUhMchD2eA8qYp/GghB/q0uFjrbxgwyc3
2VM3jgnfrD31V5V/WH50plXc2oK8tg/QK/H6iVxjp/YlPOuX1OJhZKDQbVzjw/9YZV/5JX/MWSSv
Qgk8jUyUMhv8VqrgFeeRPf8YcsQmaaTsIo4tBJKIVV27nYDaZIk9lb8p80fdRNzL0gPx6+5e/HWT
IFtc9REJ+cwYptNkxZWwWLPGNneBd4yFa3hCgsYao0bT0w80vfSEODnTXMpW71PLSlieAhpw5Upb
SjRRHZO8M8rwEj0ldTqbvEwEe9oqZ5284Wun5uvY4pIiB8cZd3DuUSWVH0s8CRIi2ctrSLNgN5OR
1P8YdYJxvnX9cQTL18V2hIw74oCFzBAa+cs8uwUZKyRvv/jiWOGDVCBo5vJYbqc71E1blanZJ7th
j0EEjqTOra72oQ0PgGtoRCkCucvdMBqPzDDdn/VlokTmVg3jmqntNRSruQfvOJ1Ef0kXm/ZY+IKe
SAXDlslQDA9xwTk4tKp/8/doRdE2lltJraiLhLfpmVGEUX8rGzXATNI4TSJ6gPsMj8/b9W97eBe7
cwmnqgqhDwwYSEmg4lvYPlGac7QGF9eKwxsxqFHbSOMvYOCJmoOPlbPqSCPbbmM3VQ3pLggtNkpF
X6TLCHVb2paFPveXQNqpb/EwVrAQKGTAQmeGPVm2Oo1rTuGmRVrYzFcfXyVCBwCGdmCZDjph0MX0
uQd5LSmaMy/V7apdi2FMtdIhIBs5Qohc7aushFiGEJi50jwWV8RmEuzA9T1xFbjo48HsXPDRCME1
cIzB0PBqGb+jxMrdsyyFDV45PsPmJjDAifog8MDaEi60lFk73ncHxT2VArnQlu8pqp7P4QXg0CEm
52AhY99m19G1s6OKK3lL3HOXTqoPrYFzRpUaSC9+VP3dUOpIsanEW5J9OHMpzCtpi19A9HMnRvx+
OqKj9m4X5HHp94lh95B+q4T/19XcYtwa/zuf/riYBIAkAh7UY0Xeh69zF3op4FO+jVjB3ZsU3aKA
slnWRHC2DriRFI/nl0TkUHAGx4Jjurgs7Gjlqz2McpYxvlKiLW0Y7QKERQd3vOGOsqGdaO/AlWua
5D6lScJd1V+5T419d51y/MNjyZW1Hyir5S2N3/sZSYC7brIaFu630zxHcXon2bl/w4Ae36mk3Rit
iN31kmcBcP1hSZ0KqeZSbPp6lEy8pCsAFELNTE8r4l5NidIwXhfplgGPQUBGhDPI7ZWEaXi5s9Ag
UrPIKn8LueZVQg2QhnssLM6tzTQGKptdENs+mHhw5Cgq6EOCNST0GSlMOJ96+rhhJD2PNoYBmIXy
HCo9kCELKCJsMJMZ8F9IK4GfjY2baQeisBF9yXg/ODJJochROZuggbfC1cpx/eoBnVHzpz/7I5gk
+BabhHvo5WIT1K+beZhXwEy0BIarW8jyShtP525fPNLlfGUNuxTj2dToEsJ1J6gH6tlLTY8q25E+
kJdqxc1zD3pLBYqCIJI77pLg1xMElFXY+kRnJjy4Qblmgmq1LIUSx4XzBk2Vp/pMohRofWjAvfh9
KOWky+vKYv+LHObMXysdb27U5swLc3/rmZy4MiCM4LloGr3S1xnMTVO5vcACqSeB6H5kN/UQdi9e
So9tNgwy2n8OGCa0H3W+er8yhTClHU0tZe2gb+2TOgvR9yaJ1tcRcIshwzJPyzaJHNyXSePAqEC3
VlzoLvo1VQpeJ3AACFVprczEcXNjXl4Ho83GWP664meV2DZl/ReBaEftgcaGzxK1rZ9WE7NR6LIn
X9YQ3icjlGy8mPnrZCSh/DcHIm98522V/RVUDzk+krnbQCMyGWe96BBcq8uatZoEgq4O3Dh+Vh82
Liu6YTsK4pFTruolKSrOAy3Nssbdbbr5Azn8Cv5En9zZZLjGUxWuQA3Qp4PvQa8GXghMSrcT0oDE
MOzJybj03m5H/gx5SEKqXHVyWs4UsySH4kvucwS0202H+luR8e2ubqtGxlI1JDmuPaM4TplNWlyK
lVrKbaCOXu2YvUnGYYWUNN/KxB4xHd8SkiLJYWsGlV4iviQRXbhhP2pGHdaBKsQ/rq+A65reL4Z8
lXkASgQzihOHDquD+QNxlSk30ZzYk53JZFmdn8OpF5b1YO5wIIqwADFXaaj8qi2aRl4RZ2RklrPG
N+sOlUDulhcoXuUHPORmEgKemwCptSwoXB5/F2w3ENVmh19oB7f+zKBvBS0/MBjbKrCiOoXKeIyB
9oLGBQABp2PY6CrTiaPCOexc3AK4QtWnAwNl7ify8OG9xcTBSflwUvy9OcBvwj0UtzEhvDqZL2/A
aL6hZdI2nbDVQi/k+2psTdcxNrNHCKQG+YV2jla9X/okU9CE5NddV4aDN7seljqTGs/PJkfj/iPa
o75HF6j8ZiVbK31RDgj3xcpWmVVFtDBTfr1xIh/lqUmemg8+kPZcHsK1RChBeDY+n+eN4n9NOLmt
RP4d3rbPT1VLK9ZOlEZIGCKotaDZfQwfm6HD1Jn9NPxFG2vNjXbb1l6lV0kNw28PyhLJmcXE+y0h
QhMlIn+l6451gdm8haGnsib/9u23QArIgxVQix/mzzG9AfHEtXLTkQTeOp88p9Q2QwA1mvJW68uc
BZtsBWFRK5PcmtdLqRg4h/g2VwUFeOeAENxA9DDGMtoaou2ceel47PLtngZb/OYcqcEzkTi16gfd
Fq01f5uerroZBYN1wgCTKtYZjMgNsiETyggxv7GUp3o6oEsxrLr3OICNATiqWcK4U2D+sBhMfkI6
hax5lsfvsrf7Ceiv7DeKUnFs9uiuBVMFe5Ul7GNzzHq1Bv3Jm9IaEqfR42VoeS/N8b9ApobWau93
KduiM5lT4GszjwJW3WzwbUEhAeOm4KUXaAuZDxSxaUK+NVfitKLxuZElrcjGBSRuEZbazOaUip3E
ibkwxuzJY3ultHP5bK4dt3pPKdYlfXiIzPqvGuOdvT3Lxayj201LWBdtq+a3StQuiHrb7Gp8E5qc
+7SxT2SRmaA41bHmrqVM4PqzNtDanwFPZ1bKSoctHHJ78O4RU4+xtecoqd6BfASNj/MgKVLXjprJ
sgFi8t5kn2zyiroHfDP2y5ToFG24BahvHR/07VYzjIyhJSJ2pwClYHNjAs70pVBxx4iLuLahxI5m
1LP7ptw4/Q6ZpNYpWKOeE9BW5wrozmpWvUB0ZoghMIodD7cVTT96u4o8Sksd/qsUQwCBoXxsL3XK
qSX2b9xeykh3vI9LvyruMDgih3ObJYRjVV3vrB7d3e3z50msWaTvyRdoie7hqu3kdSS4eTyrbWNq
qk4wgx84padL+yNnjdGoqvzrT5PyQFiUQXKdCV1YXQIcVUQfLXX0ZBHN2fnPeyjuYPdZhkUcWEAy
RgwgqSrn0CFdtN7MHL+csXqHVMug0+mPbk4zT8l7B/wFITvHZReAxCrsieOU/YKYegVJF++0CELW
xtOkOnYi1+gprfzu6dMZMN82dqzr0RG7Zr9tqi7firhCwhW3EfOc+BaBykmTmHMjKS0T/oirusvt
4DISi617YOaHmuWpM2wBH4t22w3y2vqp80siegeFBpqo9INgtimzlRl2Lc5Llwu5Mpq/9s8h8onl
EYGQdbSvvNo+eKfh0nM3sC8hz22NzDvMSSTHXj/PYsVsvGpJkuMJhgQKVEy5FF2TUTh2w7pohB3b
HIHebJ9u28v4/Pt8auCjiMzUqC6HXWxKEHNAXYuWgAC4LGy8xSqhYWyD98rz/+U93mf5vWrh0yaA
EHid5btpnmoD2MAVYvrE/Zhsw+Fw9xIuTKUBawnvCAAasuY1YGlVMor1x7kcq7477nMKRUaOJpzZ
vjH//n8zE7QrYde/LkZjAIEOGMc6UQfCIJveDOhX41msUcsTiXMIxBeRMhg8e33xq9k9OAF0XOGx
uGOqMkExcZY9aArw7wRoOjWJI/s9l2aiKC4gkZ3yiHt5r7A+ymI3KLcMhjuD2nVeh3tG29LmGpUS
IgQFzOgZSlm8bZ71fAo3JqU+gRS3rTXfjK4298AAX+fX/8SbzSHNAWKjNsM5AK0f3LDK2s9dU6l2
CtN385rXlOPWMvvxSTI/wpMopK3fcaCd5XjX9t9Sm4CHWf4ucFt1DxqL4TeQ6TiBVA1dl329Cx8e
XB1HMQXyP8/ljiraTZeRW6NkiSSoKnLiQvC2Od00tNfi+/SEC6OdGdfrur+4SKWm/TQWPYbYgmQb
fZyxvSMmzgt6mBKFeqDx6zFeqkPFLFuihRLtkWjvU1+8dUoSmbKNqD/TiFWrZh+DCRBWEVyOVEvP
b/AqvkYhI3JoFzNlX1QEH+SJtNm22V+QGDDAtOwV0v5kaFHhMpaJnP0X1oiQDS+IFJPUEkgwYtKz
QJJ5RVnkF8KX0hy/7CeoOpV5uf8WXUA9eKkkAAXjUPCjv0L/qtaict5VoWmFu3K/lXXEneaEpVgY
DS0l9s00ZswJSk9cbtLNM3mIbvdTrkwhe1VuriVv6NhC/aGmj3PdEKJLUxdYUJyCj4t+xjFuwM9m
WWqiuY9PmblXMFmDTmxmE8QD7FYap523Fi3mk+Nx/tqHSxD8tYfQqEhQ9rjpAWxWEMg6QGeNtpuA
0KqdyYg/c+8Ax3KuMlnPuIRFMaNLAeiD1yaNKXkbNq6L0hUaJROSoslunXq5YfD2RhMfoRSYqHF/
/dMIzIRjLbEUEQfmrvi9SJGGMRtZse6jZ6hg4/HtOFbVYK6We80FvA37UDWOA6ZkH04TaEwvZ0OB
+LUZ7JwU69a94KKRx6+u5hXxlhyYNDYl0xN0UZTgRG20yc0XciYvL7wJ63ojUiWPIYZKUG+V8NZ6
agshkPZ6F1MfDQpKx6e7oXfp4aFop1gPXziYVwjcSjxPdBHRGPLhSAyUkLL0pdMJBNx3j3lo8v+w
BpAgZjsTMrDwv11LP/ldEmAjkVm7xMLT9KNd01yZ4tLFHj//JUW/H7ybdsLZPdp1U0mev7o6U7/c
e6lsiIa0h0aR1CqAKtBXBUsVCxprgxtp3lZwdxVG2dqKx+SPTS9vb0GsAnwsb+l3hYPujq6Bp8TA
r5DueL+C/aWXeBrLV4wJUT5aRP+DWWet9DvnNN1L9+a362v6mbE0AZKdmPda3/Itlo6cO2Socpmk
zpcZuqBHjCiDCX/T8D1Zfo3XzMGSwZglf9Ff2mrurXmPbrKhNzkrqIywjr0tyiFmhyGHBvMLFGbU
a6yimTaO1TqJclDVBEckjP5FIBW2PyXczk03ie6ZkyKgp3z9i/LBrUTs1btxvVJBuoczGGtWLi4n
a/dDThJyGb1+hFOd+Qsk5MI9mYR+x2+OB6qYVHCAr/yqAfbb2GA8AQd+9HUX4IPQfOL36hE8+OLF
1DvQA92N1YZgHbsckmPRBxaTAaC4R3SzXDhxTCRPuGvuaqwHKO3xW+OmUG37cGrmOQZ0GwnT2W8k
N6ODbIZZrQCW1F9dAFMLzBzAwYs2CmQxUjyDreqnWAdPH/L2swmek7F/Z4nF2fbDnCOjaIK7G94V
nFYLJvkn/lMjV1zCbsnaB+Jl5103ORBnqI7ufUxVnaDDxY4sFtecHKh/n88rAANp5az3Uv9gaiIP
lsTL877a0i4RpmLppp5JW57WRd2nnT5ovW/vxUc21AopOsCxKS9F776/JgkvI1G4ArtzB7yA//Of
J7lnNnsACs2c+j2wlNABJywswM0kUT7bmVRM2nh1TkP/Hx4TNRdGr2L5wgI6srQXsK2kpJmt30Xe
UAvAQfUvAU6IalByi6rumk6otlowy7l/YSaxAWtkCajm6XDvgdXFN/tqb9vDleK5z78/Ske/4jyz
meR25ewLbogCq6cKsULc3yPcKRsh6WT2PVSrxMbFJiTMDJ6sPIwf9Nm7n5AoEarWIQXfBmzkiQXu
WDUczLPFOPBHYC6U/k49hDg7dRjh/WW7V/ksSExs+Ou4qPeghTOLmhOnUTYYz/gro7JrM7WspV3L
qKgYyG+vOJ88cXj9Au8OI5Hdq0xH4XWgMmvdSY6AG6cOsgXZpCOd9h6eDu/Yb8gCNjKKg4venLTR
2LOPZRKT4cx6wdFs0rkhQGwTHUxFX1UHQFW/aJy7YB/JE/ZQ/j/uaprDf70aPwdw2aZ5WYYD4kV9
2PSkw+odTUhvJbP/mLfVzHKLW/LYYsrG23pyPy+hC7onckqlBgPHHjEw1LisdE1qAXLKD59vmDJp
1hafbEMnA+kylfL5I1vce7oeCiwcoZhJXOd90QqcDfLb+LSTV3uz/Y1fl2bDkivJZPvca5pcZlN9
F1nESXVSL0yC4peoEEM9NFl8Nl+gOgb4Ix033ClEVWApgUHJJfjJLxdfV3nsacaw5RETYOcK8MQ/
NsWi87XyKiQxslh2gZ/HukNISUMgcLJbqpuDqzwlpFFQvKobNxIROO2JseY2MJbt1VI3LYUHFDYr
LO03tkDNCNBMFTIjnX8BTzbT90a0Sioxf/wqMKnFkp3CVy5K0Ypk2NT8l/fQOMWJqT5tm3T20/tg
JzyaznF3bUYN0f2X6yiUOXAjdNwio65SAMXcP8XiUSRQ6dsXzbZkVZiYI/iHifsYf3u7g+U2leVy
pODloj+h8SkTMFKCOUBFP85ncRZc42teQXCHwjWdQJpzRlSrnL0IybpTx+zh0FkjKp8fClwbTb/Z
884GAnG1nDloBff19sRqGD5BfgxBKPRM9W49wMkoS2Pa7Q9CRLe0MH2cu4k6vcS6203hhbRHaesG
75KBuQbLPG3wdIKL0SGZ3/BKPZqpsjFyxUZzTgswIjUc9ig/PQATxojROG3QgPfmAAj91zxqiay6
SSrVovKVm/TUSaYpGmMXWXQs1O3vkojCBHaQvmnfbAo93tPkB6wXBrRBFvb8DopXk3s9bZYdxq3j
R3yyJtf7TLccayPtpZxmbPicVJQoa6oMQXd6rMIWDsBT6CRnOhTZYDER3xhLj2cdhTKYx7yw2ETn
wxjl8GC5YovC1U9FnLWZcqLEUTDtb/HA9zgqw/8iXzW0GamKcYhGEdE+F7huX1UK9VXxAytAAFCq
qCuYI3dr0qbl8MW2rm4hZ1BDLzH66I0V6uq26LZTDIYzcof4T7xaFDxyswGZRnASNCgFSIdjnYtz
Ga+H+v4as20rQ6uBWxDKtqaupgswR0pUXU15xaLLRChIEqwjacLfSabUwgCkoTdbNbTlp3FR9ohO
TjX0dQKSmWDDfZ6KslTu/ZmWKUTOeVw/uqrVlYDNR2Xi6ou/601yfmeSBVu5iEe2Ta5y/8AWAJcc
NiWCGHk1a0Px1ej1Du476ABJhifCb7sutJTA+vsCQenm/y8THms/dREJ8n0t+tP4/wbcdhi9lQuy
36LS1NG17SnRg3joFazg/y3SHt3HgHwAsObzL1XK39sv8Yvmz1uCLXQmviQAZE+eP24AidrysFkj
fbUHYmqHyWAHfl1URtmKk5fU+ZMGkVAxvFrKch24VpvZ5ijJ74mlGomGCJrt/I28qxrkYQpny91b
S/Ug54Me1yOQ7paiVqU2cjjuWXfD5cb3ldM1hnMZbV/5zu/7KxBEdJET/Y/pco3aOBwFr+pA1SBP
lhiemXJWUJFRqwG8EKZTniJD1ZhBiqLavXY5RgKIoHulgZvaS2kwvb4fOSxgIq/jhWoIIPX22FX+
F9p9kAiDt0/OyFLQ1A6LdF8CXSm7XnMQAFM+dmX0oGfzUM6nPoe7csAStfhRnROdAPona3mMsqdW
Ocv/9IgaqbzzI09uPDbOVUWEBlXI4mBpuQ0daEafVUiy3a9csDb7MthhUwkIcbk1LbYmE6Cuno4J
dtK4Ou6emXqWR1d/3oj5k00SsHN+tP2gUhWNvZlkZQzVB6UL2hrIgx7LNN9e3Y9hZKnpH2gEtnSg
sIRf5W78/B/PO1UP5L6YMB/qacQz7ZUg43iv2ya0S5KmpmlujQHKg0fOyApWlek4y4rme4leQbHb
IyyYMc5PWkPw2z6PKX4+AYNezhASR5N6ilWfbHYLotlyS62+NdrnMBHftbi7YZBLQLqQBnCLe5vx
SYkY6Tp4siTRSjNKk9cqfifCXvSxFmxamCsEwm4gJXdmGUpRbzZl0OmExTIQzGuDuFHgloLDwudC
tuXfhO3JrQ7YHBniJMd+TJ/uDFmeLfBLWHG6das/K7ozFtwEP7icCUwYDaTQl3YxAKcK7JglFF4n
R15Y8fBwRQn0LxBMAbbwRF+8FOt9SQSE1LpsP3DBEsjnneFcsAvbNfTrlgCYjjn4UHFbRDhCRaEC
W3rMgfbOa0N/t8zD4jLTlKZ8aMmCR0+WJhmcfXpL6JwtqpjGOb2jMNWhFpuiaLFtMT0a+vuVoABj
jS2C27AJXm1C1aG6gy2dNPiB37LoU6OarLdc3yOzb/oBVA/3nJNcpeKrJVjnisXdaI13bM+lYG7S
rPW/TZfGQ6xfU7d0yO9cPNPztnLkxaX6lgktZgw6A+JWgZ/PFQrK64DyzDB1Vp0MVESdGy8Yn+LP
EPowEAG4iiQZhm88EDFbYljHk6OJhdfBmfNT1F8SWAGsKWSz7vtQpY/gBZEbWr4sI4UWgt9on6Df
wJZz/GrK8OyMmp90anLP2UWSFZDeDsN5sFYvriA8FGwRcp6YMKT/rA46fdcZZcqHh+FPRAoWKwXO
mIj4qXLPCTnkh0Ff+PodQOjvCqqgDAtDa1ah8rRsb9k/NxpE+3ZSWeinfjDnrE9NHM4pR22xrsVO
KLuydBvbW0IE7tIZe4aFVqdBqw+k52F+EWgD5GrOQXl0rYh6QY8Nrew5xD2J2UWa5rnSCU9XmNFZ
VHgGq/cVXJndQjK1YPU2EQSzV8ABUSykoDAR01tqdUVXiUGw6vOiXDI4XtmW0N6YGX+3vqo8J6a+
O8rin0QrqMXy7izaTTQi41duf8l87WwNSoKhUz9qjAvkVERhh7nur4bhsQQXmJAdLxf5vms6R4/z
vEtTZ9dOKymcd3VvUsMlvTwGYdWOXIcMFAZ5KWuwWqiyagxsIwJLlLCvn7+d5koMllaX5eSwYbMU
m+WUac3++WI4MAdNt1nsl8spakrtBsDtP5P6GPrZuoPDPHhA3B0OpEeFAxCQGfldyWX/3A7cZmd8
h6DJgxUIXty/HOc/YqjbibCNFhc5D4meAxqNwsoH+HkXifQkKTurcCmHqbhANbdlaWQ+DU5hiOKT
cBhcB2xg5zjnlCpqvMtySWFLtmUE9TpstfOoHbDUaJkFjiMyd66ODu8cS+pV5Bx3zYmtHeOCsa0g
+VKkSTrhil6v/dNg3r7Hx1gmLmfGwqDNnpPXnxkfxz/WeHDzjcu5x/5n0ihLz+q4tIa6BD3UyIdH
23HvawLltmew74yVad6AVBgum5E+8otFp8RFM5dALT/S87QvKGi5OgQIeOh1wZIr1fP942rztPWo
W+M+sAsaKaktUfm4gkxwRs7GvjJQu6gO9SO43BsSIjCgPpYOcYOnTx6WpmrUFrfvRzWfSx96z+Mi
bD0tzcbVWD1x5Ep1Smo6Z0CWZnv18XkULGuON4aQA2/S+RclJm9eWDOqr6PtVAMaXlvHiaV7d8w7
JSkC6n1yAIOVreIOpGQKYgxhJwjb1hLre1MjyWhrLiZLSQfcBR4/Hooz7IkzT4PjHUNhQHM5IyGz
GFZGQTYiTsD6aXS2sEXqScCbuAI9IZuoRKVVtPaxZVLoJxTyBs9LHmIStxfkhkgxZYsOdP9tjtl6
MwNR3uVhBL4nkyu7nlNb8AMVavtJf6A6huA7ysDn+sjYKiEscw1LLx4pHTQOj9BjmoZcG9QsDjhk
CTiOa9cfwbMHlAnQOAHkKn6CAhL8eF2hz4rVdaDcfQxuEffTEj8zTJjunuiCWYFGln43LaaMXtb7
pNoBWYcUA0WxuzyqrOF1k15PRXmbwPK9WLP4GJc77SKbXgktdXiYf9zCnsWyKSO7IHphirFALHuc
pJBnp2nA4un/bkHTEEx3ILhEVoazQDMwcRqgTjaW/J6okJIsUVC6YxNCj84pEfHcJngtNrCcZzW+
a2NVz+DSqiRE1akUJ0WDdKY0V1vCifM8cHOsOyerhHx491C0L23a115j7QZJNF32Nht86fvkdUj3
a0V3NryfhEjBPjt0p91nZX4NQwK/da2FcR4GNBgNNRaIo4q2x1r5yf9i/XuCkFyP/PP9lzgwsWqB
FMzyWBiU+3xqVcdyezalrRsgWALHDfspPNAMTU6LmAtP9zFHTStUD4del1Dj5aH2albJSYq+9haC
+4w4GbCCh0yzrDx0AeQ9YumXddDFqSdsbidVI/XEjD28q9mZ40AXNkBpxpBdsRCt8rvWO5ahq3lg
pkr/+Rp3bqwjBMUPPYcrZJ6SRkG3iK4xNxaSXueJv6P3GqUAtDWSGs0q7PpTadSWUuoWdwijBiOs
E/JCmq+Z/WJwxb9DycHHYUT9JKblO9nK3x9GcRf8LTkLEJ6RNPL7NMaXFJ731gPooqdoPulqV/KT
k72k0nIuA3gjSN8b5Jr0DN0Ls8DluNqkM+sowTWKackJtBEVwb2ZsHyZ+84ymf1XL1A7EEHYZyhR
kk3iDFlZsie4bZq5mZmyrSu7TOBZgEkEFr4UTwJdWiHGm2oNbfvB7ujXQ6XYusRHku7IPpNMKozf
8LsUd3AmxWWSy9B9oigqyNqL2meJkYOJp0HivV9fvkVCfi0cXLlJ45ds0PWXOUcNbye6+qF3xZTr
Yw/n3WVubdz5xmWliLWjhBwr156qvqzWkiF6Sg3L1y/2x8VpFM+GISoXdRARKQtmkT57Rn0WmVA2
GJSZHTt7ptbkUfRxW0Tgp7kP53wdnoMLMQ9Zw+/O15CyhqQ6vAQxufL6GKDCCJlq/l4fuvuQ/JRx
HXUvcey8AoTlMGjzQNxwLbEOZ/XUSQW/ugLUJaxKaTsvUmTB894qUp6z9FSjvaXBH9CS523ughRz
ooRbUAlPTENkYvTdk2CH1Mbivkxd1BSWeYjiQKJ8J0Yv1Wt6ljV6gmEpAFzucLgJ8AQzwyGg7319
lRpsvDmG5le3mrO/1ColzIs+kSDOVJYm+98tS0OY8s0EEfGeVcwdF7OyV9nkEIM5ngXW5J9uwnSw
Qa66JWyv9dsyo166nodZokbHaRZ9mTYRqknsn7tjfkaLXLB3ASGtchanmEc/s1BcbzXexxrkLQ6n
SyC+wJJ98XS38WDTuGLVcmQBXd0W3Aeu4KC0AXnv/KIoLD8TMbtHzxDAy5324D5T53MlfNP3FEMC
mxWcWZl8oIxM+IwlWMLn126iNMFExKivdsN56ih93/60GiigOzvwF+O8rWUYJ/BqocCvApiWV22z
LGLQ/DcOD1xyoNYbqCNtYbcYP2rfE2pp2ChgqHH1D+FNc3h8t/+D2vI0wyx20eqE5Ic2/lVOIwW1
SUohdY/rCWZ4XFJyoPn15Sjt23KIJ/j9qyf7/oxG/U2IQ0ZZpRGnNhWjBP3DXY9rlHFHS3TeM1HJ
reU10zvereGRfiaM1HinsFuyIDDNUfmnqYxPHhWOKznU61RL27F1Q9OLzpK1JoA/vQnfb2tGW3FN
znR44Mm/cXLZKJoKZw41Olqip+KXpvw1zDEPymIC+wIrUHqR4pUyYSDX2VAZeTOs5IUZpb6ch+Q3
bEqh6tbFidwT9QFvb3nkouPlqlPXw2cDarq0FV99xhA8NmG464QJHHBqEzwciSNi3Oi/cIRLCUsz
x/SdZmUcrn3WAUN/gBD38NTyu2wBrBL1wRCblKsfFpcfMvnevnl+wzAsOT/B2bK0BnCFNQKUG1LW
q9uMqkP120kAa2mzGSnIdy+G9KfstDZor3SP2iFOoLOae/XzHDh73qgAvi4AET1I7tf4MyZXyBpO
0oFeFyx+MRP98uyJFkulj3vuPT7VO3+bSRtxhPDotRu9n14yfDgGbfPiGVReM1FHVEB6Iv0+tqDn
Np1GaBhAiXGJIYzxtR7WxuiXDve4j5Ms6F/F/ZAtde9B8D+6LgxKN7zlzGmBJt7QgvX85jHKvAzf
x4zdjNb8Lsjxc7NJaZA8Ok2PfJhWgOx2RY7IOR5UJqI3wuQ5CXnB/90oLDbF6g2ATbqej0O5DIDM
kFg6HBZiHh9OTaBitmGYS3JscpP7CCOOxgnS6/fkEBpXUbz5az3ciXhqv6DBWjBqDUvJLv5qEZzC
X+xnUBXKOzY6//xbNabnsegmkZgnhlVTVOVOrR8ow43IeW/vCzWJ+MjpajbzrM4H5wdYhZ7wQuCj
bLl7M9hSAFQ5ch0aHHpv5EPDlzfrZhAscikXh8CGGFScjXwNCfklyZXTM7fBoq5qYhLsjnWDfelh
CBC5kO6bdCwjNTrmci/tUafj+ASB8boT+Nmq9MZ0DvmcuTl+2bqnKXyyWLrlsXLTDxC43y7KV6Jr
o++7rmEzGqFiUecot1c+qXROtP55hYK9cfyXfwSdzU1p0RXTCq/04bPw0fMwiCv7URZb8aPYYdWD
DZNJZbwAStJKqpuOTiGFVtSFcivDtpQE5DlPdWwWhoJWQPv0R9VESoeqYWHr6h6GMRuBOeHPf6Fx
JLeY7B3dkL2aNSrQ6XxENfuv6x7zaTbHC6++1h8Idbe8m7yOzq5Hu6DnHkDrfz2IyPXqfO6E+Y3c
CQFiP+CYgLQwdlX3BDt/gfiKkX8VNqgSHl0daMJb8LC1Cg/yv5QftmadG2aiM0Hyd0Erh6BZPJ3a
QTqW/qzPyZfjXdVuEnvLIFuABmyd0cr1rYimUWpELSk2uq4gGWc00ayJF0rvIKfaT4+zKuk7YJd9
Z67uk/kM7WJrTueIeWkEDREA4JgKw57uhWTLjnLExw366UD9D7UgjkLfDm9ibWAbJJDUrLMzml7M
WANh0blHK0YNkzDoQlbkbW+MI7yiLl6T+0+VYE8lmIRzLsAP4fY8McLqccnKlYruNwS4jjfY0kMt
YazJcMNQMb0ngXkpRLb+wue4uoNdGv03uY2NAozrA8rWA3VW6GkMaN3lpZvnAZNR/eCYiWrf1FxP
1DyFZ8mdV1JgFGOPMbXzxRqz0m0LBWoYMhkTAwQctE7isvv2fENQRD6QO2zYrHpCRAjUA89PK/RV
Gtdsl1LAJUkqdK1/0GQa7E8jInqOKeQAS5ATBJVljp9BPVaZuf4LTGaBW43cIDdxgh6tKgrgpiDg
/VMxkYWzhvDxBla8RvFSbqlNIvJN12sZjp2vkBjtYGbar72wjZC1EqDsNF1OomkyJ2+YChIHgZi4
lhmhpSG12V72M6w0BqbjD8gG2/FfQEPQfInE3atQ1/WMSQf9M+/lx+jfxo9xIhiIjK7AyOG+uJdu
GS9zDifdT6Vrywg2SzuxinedgXfM32eI+1efY6Z2nxP+EtJ2FuUXrjPenX9+XWVatQhrWmXrbxCH
zvcwqO/74mpcpx2snuBVCab3g1WpU3sRe3EcRlVT69jzUcCuTcDonUrBPRbIepVjfOBucbTEFpcA
rsl5TUMkPAHe2zYFJlvckBnAR0oLdLYAbnBEwjQWtxxpk6Um7swYPHcrX5ih9vIl2FcKbS0Lpuf/
RCp6dNjJ7fmhDbIfQcCxBQF+h7WZbPf0l8c1D/iz25NDj5zkdVcLkj4iMVxmJ1tRGPKtRexNMal7
5jHjXIolTdVF8YELgdNJ/dN4hwQ2/s3fuXjluq+Qa7VfPqL7MZDm5H5MYs2MHv9jvkTbssXo0uMO
zSqsedRfxIGzSl6dJ1GTjj7B7gYWWlbIEbtv1uPv5oqKanMcb7R5V6jrM5e3vmroTXm7RnxS6JiX
q+LaVN2tg/sygpxXDqbEvVB2RnDQAsvp+SWVPgnRB1lBrGSB7LwWjsTOszN1fSLs4sXD6a072L0/
tP2EXOI4sGy8ZATQx6I5d96RPHjCXoU+Xd/uBsKIOdLmtx5uV/qnOZoT0tOAd1WRBuA7o3B1Pt3Z
gc4/9j6ccJC+tkSSqJFZ/BInaZSkW5Qnj+xWw5wA+FCAYkU5Dik2mAQ46FrotpEVGoQ+joXyVz1L
e3Snd2xehifk9i0auwCJwnBhxDtVcPAydf7fq8KKUiW5jfo7JH+SKy+WfsczyDYckkEdfrFlxRqE
6ypZYatjjPdjkkajAYh+XixJS/aox/tk4IJkbqAsV0BDQxl3GI5mOGs1maMzIZWEVZiOFhH9CMOO
QZr8He5iTClUstgR8kj04+CM5Y9ShH+IckR4OCTGGgYGWLXRM6OrLa3s50C/JTtaWKkYhox1YPSb
r/IIyfsyh0v2BKA00N8y32UFP2mdCPWT7+82gIodmXeZCAqQTbPpinccpLOcz2jrEyAiQHy/Xw3F
LizHz/8kT8M5mFBmgXsQIgU9pBavNptwWtprRV68raeGT9Pp3yVGkXGSpYnH5VFj2fRQlHPjQtuL
nkVgA0EauT4D3DiW9niMnQSxDHo0hLA2tiOuC88KG9HAtekkl4fbHA8m3lUDFqvkIv0/+oUO/Ms2
BZPf5nbX1YDZIl4oJFLnmSpFyc0BMKByTTTGEKDcCGqUISkJ/rRm4EMZwpDhC71DVfN77dz4TcT5
DiY0H/bEFDJ3fzP8g89DW0amc5LHf1zctUPf6coif+77nQp8lP3uMhDT3bdDMI2Vkr6Q9o6ujSc7
RUHrT9f0ujGrMHtlK9S/RVwZFxIMy14bM2fbSVlPsBqmz2IIWZiMAuJkLELRE7HhVns0sSacU3Cw
Iz8auWqzaRJrVVYrblTo04vk+KHimrtShJ8FagGZcZ4UQqAmO8IkO+GC/lqIQNT00B7RIMo+6fGk
ktK5NlcfsiVR9iHp+sS7QOk8UA/7QXxStSurVykpoRPS4SLNVs+2RQbJJ/91rLb0G/r1yrqqIDS0
dSlu/JVoS1/MiRKWxHiC60UMq323TeD7bZJkHTGv6B1em5/cO9RvuEExhdfNx8iZBMmW7IzRFpP3
BtlTJkkIHXxOJJIzrLWQ+lvkOk2c2/UGgqdQWd0Mb4Qv+CpvRv8gANuFG8NzQ+Fvmc/GXv4O3T5E
cbI/Bd+suaot/aJF3nNiTkapl8XQ00Fb3ThtmKRMTtP5xvzJL+h1tRkj9cNites76bmRi2fMLAeZ
0+0tG/R1gqrs8ZGjkKa552ZrsJ79bGFg3cur+OdgtMBJbbwdgjegPNV/GBzS2Ob82IjZDYETbN7Y
yMNHwFQnVEiY5uWGitDU03/rEFzI/W82/sDPDKtl+JaxBR/7rkPX1tRaiBQImGcR2btr27tXy6nA
5Eu9XnW7tA+SD1UePXH+VLzvmtLm/6CTDd+DVnkUCaEuy91kWNYqr7p0fx3/zUJ0HG/Ud6yGma4s
RqJ4Egw6CpSzXJ/j6N6imnNJycNaEf9MC2a8xcq9B5apJK0SqVbqIPOBLZXjAqu+t57d9vhWxtti
0Quc/PUoDIM3UUtFFrVImTJNaP8uxRUkIzv+rExjfXH9FJBfhhAWlWJRD2rjI5S6m+HZzkeQeYag
a6KMwzyOOsVwEoUfBTHYVEI6nDffRFPOyiijIhr1m5NXFGZROIhghechb2N3RpblcYI23/LzjpR5
SPhTHxd5aduMeYX5oQZYoDxvVjRBb3uAHO+hP840PVeMuMFVQ9BNYA07aeNsauNMCEwFpQREk6o+
vEd/J25czZcCZKx3f3c5kjzEuLEbxLlrkavQrkNELaWJl/XjNFUzK4X7ArLXakgL2B/gnjxWoz+H
ReqhVSb2eAfhhcLNV3OZFOdkYAhFpqmkRzuYgTxJ3TFu7Uoazpy6cHNFGlsqJGBpVuTvYCiMUWRL
JOSURdJX2SqE8z96jPj9ofwsz5prrc3FaabVSTT+eJuecBz8UWn1RiP7Goe57xiPvjWNhHpSMYnN
QZ3zEfHDnK1gqsVov+G1rB7+JftPTKd0QkaCQH7azhqxlLfBxNNKID6CWJwwWdWxXEVg+NRsyKHJ
YeC7oIEQ5ZIR5u3eXpx/KlMKZsdxCLJ1ynEbC5riKG8DXVy3sZUlXHiTEauPkoogao//rnJcv3iW
T8CApYy0NLds/UWIQYlc1EBBB+f5GgnjVx6sKYRhBzHGZnXTf17EPWv5zdjLVm1N4Fbo/2DKg5rk
km0r81v5fUyFiYdIi7Tuc/rzqzT8BuvTIo7k1YA5D1Vn87gcs8NPOFGObyXLGEPV0wHOTAOeNyuw
KuQUWOt+lfPhDKE+lChLjZ0ge64Oy73J+PdvFQtqzgXdNHPk5LovQ/tc9HBYcUrZK2hnewwfGqyl
WCp+vLy9HwQSNDAJAzFzeBR9mS5TxfPmvIsgZyFdntYXE1X449AYsHnJg50kUitlAUqUFxSnpe0I
JszJ08+LDBOlb539n0e211r1uHfm1KoDxwVqmY3se57n9GdyCLrRN37w9f8x498jXPg1jyhOHDpZ
V4uJmhrgp9tT8sWYTTt6Q7oKi0KLfUYd6MRm2ANnd3FsT4cVcLnYRosllOgG2jgV14Cvs4f/gFS8
fHqeo+LbU1WGgUCFiNgYxJTMaf/8Iwc7em/J2OqxXwk5D4+Yr4uEMdnohqx01WyJ1G1pjX1lixGv
jbuertYNVdW8vmIPS056bnJIFmnIVzjSg31XEKcXM5ym2zMKNnvviPgdKOzJhQSSfl+pCTO9OG+u
FOZYM+Qk3FSK0LZQZnLL8QnVunz86cRo5QO8arrExcHPunQAl/YTNd5bVYYTLCCz7yF9IxXyMih+
hEGixN+1eai7VW9V2OWZRL3I6Jo9MucE8zMNVIZAK5/rBP6kEiQl9/SlXfrPK+EkfGa6ZbTq4yCB
2Q6y6C+SUl4OT+d4sfSQioHV9Xz2dWd1qsJ8mLfxEanpncnEeL7Mw//yAnNHbEH/LxuDRs4YJxzt
7AMLDFAqDg+LEqJ9wynDxXQezr25Vk4tIuNr7QRC1B0FAarIQYwA1ZW8s3FFM00Q2GabTBqH64dm
9PgNDpm3Qx9ndCOQVOtCDkUYQSOGDAPT+sFHE79Q85cfCqE+b95rt2ytvjwVB9i9FZJmCWuAjch5
N2TYb+IGBLvudoDDo2P+msqRwVa/AAmwoALe26TpNXg33KN+XFNnmXxTCJbPj+lTHGf665Nn6wSQ
m3XFgWghBM51jbjti+EBPodDf3SZACu3x5cyGmguy7eFOCtG0eX6sz6DjHH4sER/r3dPNEtJywlN
XPbDWulSNwwhu6yMwrpuIJdF8avsz2/+uDm5PbJCphrJKYLtYAuxRkgqr4R0Yv4u/z9ysuitgNXC
UXz1jN7HO5js4nUcX/mbj03C5dj6F4b/tb38KOigz1DoBFy2ZGdxJRm9ceqEmDxwsmMj6FmQATax
EPqQIumhDEtct21NmFQDCr/+NvD+yYR9ypa13IYHzK3l9Tlq9j3i6hShk0pC977xx+mxxSWg540O
clyGy302kvG7YJkNYpipF+hEfyZb2qQwpaoGY7VOZ31tvLJHtGvZMjkdM9oDracF3aC0ygqCJT2g
6w+hA0n6ZOQTKQRmjKAwwnYZ/sz7htrNN0OKxEJcHfZLWOJHpLx03HMbrmq3Xyfwyva95IkRS/ea
MvtuTbFG+ffKDHl9s61KYaTg9O5DlZuts7GEwzHcM2nguuVS1WUbDQaJm/TTdrRnAybNx4qkOq2p
ljtY/xdOS2iJfnf9BD5sTr/MPVsS3KaXYpfnn/dFPOGIpKC6ys0IfFQibAg6kIkhpweUFbX2L+48
kj9WvwZWEsOn0E8NAEn95JWNRVP7l+tqfkcGfCjuSYkrqFi8VsuWYnISP04HBhiCzzBtmEEeSC5+
fSTrN4neCEw3Wenz27IhQeLc15JAWOB0UyfnWgfr80fO3cWxfqFrNZR8z0Zr58ojs/8ClQGbkbNi
/I2GLcg3Qu7DB1tYd9FdLDAyZ7ktqZFa+PMGe5v4Jcml2HEzVKWPfOzzxzeMVlaCrxgSgpCxovQP
Q8k49R9ukRKbJU66SSOyNb1QC4jyCL+Pn1TzMQ46nVedzNUZjav0fnUCVFnNw1tRsLJbIJlRa5i+
MoOUMW9B/y8s0ApjiCA8sHoMD3Ay5QW/UpUbqm5aIf2hwD3sUS6wHQhdq7BY7P1vSe5gkkzfnK5l
qHZwpH1My9s97tN31+/Rdsu5yefdia1b1JeF1tdqtFvOK1FpPpZz2hkmbj8Cs03Gii4emG26TPhg
bmqEhD+Bmi2t/xhgSf1JZ2zs6vmWJ4m1i9UzHK3gwEaf/SZxgCSYvlMWZvI0sW/py6eJBsnCfH5K
sJILy7UPTELR9x7giuHcmm2p85lHXuzUnX944ZsHB38/S+rlN8hF2Iwk/wQ0j5graYkgsH4ctXBD
m9g5/aP6on0mP4w1tLoeIsp/+gArh5wg0fXz0dWTAkPGKSClvGvBvlfFx7e8TtC4hWtLSuKazZHC
IudUmzIPhx73tMzdT4GZ4Ot0Hu0sOZNNadL64cDcuKkj+FxsB2xCpFfPLShq0J2/+MO3udWT4Oy1
z83rzoGUSGinmQkMn+H27uCacpIq94iVGRDjpibfzPhLjvjeTCNDEco1J9iWx2k0xwt9kinRKEwp
XPmDrY715DeUb5pAnHGGy4RdMaAlEzXqrkfSo7O85CAsu69meMbnv4v1F4S0CDD82j/fKA4Pd7XO
rrVfqPxTjZRIwBrnlACXaf3zrJYvVBSSfa/UJIfyetMReoHCfiXu6kqUWXEa5Oh8QWi+/ecIpmgw
R/uQiN3OVNC9pcuMuVtQ7RyXNmTvsZovFRDoeHbFD/zSHu7Er/ADXRDdMBV/i2dd0lXiPv9mLNaE
YaXuD86mvh6WXURhsYtcE6fJMb6t5f3mDrG+LOq62bYVFDWlGDn6WuNOY6o0wdY39ViWoVH/iG+7
bDYIV07ffTlrBKYSahIMd1zYSMG+tOjyOWjQ34CirdDbJMGv4SXsH7vq8bGXznofGUheLjuNfINz
FJiUFGlaos8IyYn8+CQ2ldxeCP+0ujdE11+9yJnx39rRL/YXaCDexokfIuzRBkBnmh2QyTXuqPZv
EpqaaljjNW2Hw2e3cWkzMg9aChFjPhRFX7+uFUTBEwhrTjlxqid0+Lp5PiQi1XTzeGxp8+5VBHsr
R7+3b7fdLDk2qGwLVXiwgu4IjtpHjZ6ymZnPaDcrO3SX26GMecj+10+vn2VBn7nRC0Um44vwVakq
KtGZNeuirBMbwPi2smsZVOLx8ttlBqh1VWFkbyyqfXCKQaJa039PdPHC4Bu1qJuYsdR3+ciz2L3s
NJWQ/CvLst9gpn7FkKKCdbw3REjd+tgMbmgWg8DR+AScLPumMRYpnQk9697uHVIpo0X7aRlM7nN/
X0K/ERy/Y659ttlnUFM972Z2K+fKJugGW1OF2nxfR3wnPFm1rQGd8Q9Ucxb+BXz2IYrB3dPM8BPK
Kn/FM+QK2HkhrzAiUPEF911QNR9lg6byNCsagjCEKaTfzJ3vTqL6jXK+ZcD5TypW0J5ai1lqv9e+
/tTuzRFbDwvD77h71YKFxgPJKFxQc6YKfyYrUTpJoQM13/5stIfY2x/Y8oPyKZhDPIeQ5NZIzhq2
Ex60bnBqZoTns5h1+sH53zXmG2UOWokZlk6hksfJ8LP7OSFBdh4E+CI7qqvojdWVEG/kyZeJN6nh
BiVsoo7BLe98RcuxXJ/WF/VJSQ82GYIfDhde8YRSNY/r7TDyCsD0AzPj3YFqJ7BIGwjsY4b41NUr
cab1x2Xxl94WyJVi6bFMTFSoP3SxSh+bsy+pvMTd3LGwc3DKKKrpjPkOsSqq8Z5O2CE44PujLpP+
Ax4YaKFtgDC+IeqWzDVmhyUxC4t+T7lTvl6AwoIriToA7kmmmBdxkdVavBFhWv5he2qEOPuTKuXx
lP8lafPu6sSA30/3Q/enlZqD4VrPOWQWbBSpFdNBkht56lmhiSObP36K3Uy6W/avgHOWeB+5hLF8
0aVL8BaGfe/seOlbFdnHk8JoazgZdml2G6SPUsBVbvOP7hTOXWOSyT+3FeG1TpiOO/Oi6gaXrJb0
ikzj9PNrx0iQgAVZ4bPMRJnIN8pthZqhR3NYOyrK/Qz+JEPwD0C/9wfG5OTN1MQYKrG6RO88FuXq
ksAfD0D0BH1rk1lLYwkWy1BFWEyZ8MlJq733Io0N7iJz1h9rMnsKil5TDPz0hkszIdxMOhJBh1fx
KMAZKSyUQPEUqYE9mxyvNZSt5S/JYehuFu3mIw34XiLIQD+kW3GEpv1K7tXRi4zt1hWbqZjwY8W4
du55Q1gSbYEGdnsUDIqOmYgA13AJbwkN4jeoBJrSaMToFcylr92UuZhnzG+ixcb6CTG8igLcNfyY
T/w7unHXkgdE/Tu8VtgIfMmI/aQCIW/IwoU08WhtjvAZ38Q3FkjH8UOOaCVuOhEFYYd8johIz54m
ZAgn4OoBcJMRJIMw18uZ4mG5Mg26WGbI5lfnenDPQsUbNm2FsuJIb7Nw8JpmP8NKuupkJIMEcLtM
BmCbHnsBtzsV9YuEbmEAIJ7aJbRCPMBGKfYZ2nWHGWJxEAVpZZ4WbPOlvGI7C6mkfG+RPYMYea8P
XtZg8VKDOnI0IN/dhBQcv2IVgV8xlkg1o7fJOHYC/4YX+zMElfHkyaV2yLvhaJUAGXfX9hTXL/9h
x7ximAR+Qo3NhqeCY0VEB2vfLJ6EWih9qSRAweJ8uB4ZUIxDktVdVETbxeX1ngY7Zhx0JdABiHEW
SW3c3valWHg+aKaxT4Ei9Hjn+0Iny5VWAsHjW1H0PTV6pK2y7oAu41ghqLlsKa5/EhBp3AcGp9YZ
/9GwMxDXGdkTnxlBdKCUoD6vHuqvYBmo2VX43BzxCXJ6opmWDfroyeL6paXv+z7to6WGO0bKLU55
Q+07ysjAaKR7Hifv35VDnk8rbifZdG+cVLqoo+FtkqMS6h3DF2LB3MBkuYpDE/ALktYvhfOXdCV9
MhBwtiZt+9fc8LTStUnHq/VcSLggKcfWZW27lzw6pzKcT7V4VB/PZW3ja/zcHCaG7xvfw/IFnanN
YSqBSNJeYDJKiPcpys0JUrUcpT5jwEZb4gJHgZxpRXdlbPKroK0l4+ji3LsiMQzt9U0mTsY6TdA7
OqKOziidQqoS1nMS5NLlpjdQC7I45DNlTIZ8gOQojoBzk4iS+Ra3c9I+HSfkRQUz7kMC4eQzcM3/
rQdfxi8F5V8dQL81Nyn0uM5iOSMssp067XopKfC3+6GRBnqhpRSOoFO+UshGOybk9+pe5R76onoo
Hyyr/HTZzCTZV1qf6jAEZkZVbZMOgDmAZhHeV2Iv0L3YAUSKJFB9XgYwC+Z8KbE/eodLJZN5tBhR
wpb2Xj46dnXh40a5LiL8qqHgAJF4bd4VnMnEOZsJW2uTvBoHBChOfiq6ATUuE6c0jfhCz4jlu/Kk
hnSQgzz8NigV4FkI14VI8/RNEaJjlOj76OCip2sU3ttStVYwlMxR587SZbRnuvJxo8zXTTOK8q3+
t/g8rhsM8CWBagQWzqHVDgp8nnVD2Ly+9w/RjwT9BFWRQ8Ke8PdIIZt2lCpisBVGJK9h+HoYNIG+
zufC6Lv0HVlopOd3Ynzi3h2IrXSy5XhuFDjz2V/2qaXTnIC2N88Bo4FB3P9uDZ55P/yHixkpWL+A
5HkIV/FlfxJqkNUbDf6Fn9E2VdvQYPPKeOQidpLL+hnVykoEIjauBKnmi8kCvK6JbXttNtnFf5bF
Pw/pStlMF4SXJ3XW4D0pCT0ilTnIARWjP32V/PDtES6VxZRqHLifgjl95+j5x4OW3P5x5kG2Pwrj
iD7NXiQ2ZoIBWP0asThBpWmiNfGq+mWjsE722oEyyHLf03odv6H7MEXMlNrW8O15/ob7JxbmuxDv
HP9WWPooHTNCzpCTk05WjHrid3nVacB5mZJ2RvjkAcxbUyjUnA2um0M59tqHnWfTarSNQGQx+6vr
36LXjNK55guMlEnd4ZbluVzExas9kuYJXwadbj1IuAVbJdBaMkSkp/ed8ktXKGwPlAoW6VSfynY/
XBfszqa6Ut5Vx2Wm7E0zmRdak/kk5HToMH9HVfZEzBlZN4o3oQkWhCTsW69pjwbdrBu4ptBDVRUm
cT8N3QolLoFy3Qj+4OdytWK0bKM0A7+E5Rb2Iv4RQqVSb8P30gmeAEc5iReHCNkkW8kTXZY73AhV
tPUq/gDiaonHLHS8NyprjQHSjVtjTSEyTmGsOTUhP+vMS/fsBD3jdSyu792mqSdEUXICmcZA7+PB
A54LF4PKzO5gQhhilfGqJ+uRHB/HsLkKPT2LrVPcUvhnDIB3SnxrKLIe1L8DsA1cUjhgty/0yBIm
//PQiUNLqh9khmIwdQzG9CqGYqotCs/NpT8PLeBbeX7Q9Exer8e5g2q/EnlTCmNzSXwadn7KGPV3
Qxgh+Ms/mvflNpLJhx279rRt7QE4WyEisg+DLz9yzErjxw38Z8+qpVuDq6JOzbfJfiqh9R99TqHj
bEdXSSo/o5H/VUKIhCO1StflYUZwYh9XfSK6YQhDMp/BlynavzrJdLyhNFRqWiYJWIxNEfK0OxTr
TYDoPZ//WMT+BpMy4mdrzIUt5eDZJ8ycPH6iFL9CzoY7bOMenvRBps6mZltwMvbb+iwG2OAgaH5A
eU1oW8qFhcpAGPNNNT7cvcB39UsG5C3Ijr9GWaSxB3N0cpNEcA+LJHjanO5omePKySubDNYDZCqQ
AHrMlixtXZ01GZPxK92SX62LDtX2QCKrIgWoiPHfsuxUwWjnlCMIdVIzmo0vt3zGJKj60saWQiZV
7+eIeNdwFhHyhDcVKW6ThIBWZ5ZA3EjWUMBPV8g94Vh5bRsqr/2NQvwIkW31WLiYJSr5+gKLqDiW
e1kp+k3yHFvzjqxRFbKnEuo1TAzFQ8QCuxsJ+jyFR1bBVlHEQUnpV+1G2AKIR3B9t99CwZ8QFWG4
sIYBgkp0ZD5C3k0/0WRT1WOVxxjmV3/ed40Mdyyib0IfR5bxgsRl57y7ye1t5t7/yKQpyWzV5lst
/zRGfG9/PRc4Xb5nQ6MF3Ld0nKfEhS/fFboXGOBVYwe1tPpHM3mohu8t9niAk+98w94HH52ZtRcn
UnacwOqA/ookY6tglImjGqWmkrkfK+20yesvVXP6kc8nHPi5TqfyyibPP+ZmSTEHwGevHSy9iyoK
cDam2dJAp5IR2PYb7V3zUmFISfijJWu9/se2P1+bcIavsZVBLCDi3lvdoQ50ZSp90kZfD6Gf7Z+d
5Azi1kRy/mO7JbBvHPRC1m7zoU25tDSE6a8lQc5X/L9gtjnTcPtoMblMqYHIevk5z9QF2CLtNNQJ
2X29f4jJCrAlVQTHmE6XxI6V82klKqp0fZ2xMVHBCWYIB2CV5si6AKkSlQKHuxd1fWMdShZ3FZD2
EJGYua0Of0B676scgIt5Z1rgQL47p7BG8zhHNpai/YpFuNk5c5y1b6UbqBtwpOvKE/kT8twTajSo
pJCmwX+IV8KevDH6voQUpCg2Wy+VOpwgLIBBCBrg7GXWuAv4iYib884RkYHPXtKU1Qgutz8Xmb62
0qLCZxoN+Mb0NWvAqnipqa/CaeR/TK3DlYpX1RxNZlKtHdopznZwVp3gKuE9fNHfzRIIC/Bwb6pe
TDtA3WMrHRlXV8G67Z3N8txTSVSab1bsCfjyUdP4R0VUVtw2i1/Q6ldVURObqHV7zmIHpsPClRK4
txNGXL7L8LvPTx0VJysgFGGjVLDIBk73RVf0O8Qbj5Cb2tw3zHXVIsIbqjMRZq5oNOH2fT8lBZJm
WrrngXi+gByrhS/1Zk9wWwvkvbgfohVxQYeilXMk44IbPMPGxS/usSXLG5oTvI2k2tuj+rAG2vWX
d8v68AanF98HP6SndHbdHCrJKfxTV9Y6weZNVUAxhOkqrJY7lolEV35VtvQ5N9Gzj8LTx7Jl61F4
v6a91NolumN3DqjHfPO7QI57USQ7Jy6zddWswGNPunZ2xeEJjTyNkuWw1aqLOC/0Fr5q+PXnth7k
2MR6F5LwlM4v+gGfYKwLxNr7a2KjmV3XjTeeAfvrdM6g+Judkquxq110UJJzLVKJ4ryC3dfXUO1/
vE+ol+1wrequ9OVFRdkHtAzHWnGjarZZpwmofiB3pBeGSebdHji6E/BW5Exfk5Lzj92ZSrJlL6Yr
UI34ho9qZVUZQgyQuLBtYaezwWzdAFmIPCheDGkH+H9X6mBFBJBi2pkvvGpEvV7I+DK1iiNlcAmk
2W45zzvHzQYUDErJWesyiV1+XIwCuvnzsufQ8Wy5Y35VyAOGhZXw1SgFM3nu1v3rLvt6v+v13/rJ
lMWU05gMV7TAo2Dieq7rdULJmI4dBAO71nxLd09YGDFiFFqWO+l6DNrxNulLGPVDyHO2MpgKtw7H
G093snwVYdu9M1GX95XLOxDLKxtcIWy6cuKpESF2nrQZqEdF0mYoOmYnRbZ29fTIxUGVqfbHtT8n
5fMFl9UiyEEl4tlEhkoonFHfAxCZd07v+1I7nSqSlEF5t+O6DuslnJInzLJzmYwI2qhyQFc/BWxk
hCaP0s58TSRjvI3AH8/uab4YEF5WQ6exW4NhjbSqNxFwLuCoff6jol0uk5og2qQIuczzO9URleaP
Owpg2bUSrQXquYx9PcQdXv68xm6t1yWwBGYx5f/9by1qcu5J0kH93NAVfUvHLy1xKKF/13ttcgUS
8jT0ofoKqfh1ZbuTIVvJzbKJE9cXdfvcvfrTBmzXGdRWyDbmJhiSDUrd8ZKjzFahSbFvv2fZUxG5
H7OpOStniKL3pwPXUKRX5JDCCuxPJWNg5LB2l1AckZ4wH2SBwKlRVWEM71aRe8u1ZQFof97O3GQy
BJwE2EunkXCtOFD6+oWyJiEjMDY4fq8gyviXn0zqbGw/5Kiahyjr3qB2l4I6syJH4T/kQ32Dj1Wk
lo0zXJXW/KWbS7xBgOxF4Yqn0ApHBtR9mDLNBP64og8MUXpzjpt2cGnG3Ei9jqo5TFO+WWWPM6jB
PdkW5kAJk2sTznYHgqJr5Cqv4H0zOBiStMeCKMMAqC3BA9sYGinkZKWysm+qsvxFyJ0CiiYcx/ts
swC36fX5bXgbf835A6Ph00xty2kdC+PIeZi8pEl4XLPt/DScpSjpq6szM9EDZdo0FnY1k0zDE6Es
KMFeL5ghpbrtsGSegwpE4xnC+zSJmHmc69Va7ncnkbovSnxwfRNVrF6QBamWLzCydjCviWa0S17/
Kr07XxVl4JMjM70shC5mYNvdpAcxOCJaTgqEssvU82bndDiEr63rKqSwzUO5a7mu4I6ZljOnxwsi
zBIMg41e9z5BcriaUpofc9vGXmCKC1TU6ViY6kQHxjcNxbhETf2+DAeeSJfXsiuW3/MyogqGBq8a
OiZr1R89k7pnyLGVt2QWZ0wfFGMGyncmgK+C15z5tpMkHqcO1v6vtQnxAIYqr/qwM2tx8c/+fa0H
tPqKW/3cmlWSl4TjdqmafZd0vYUIPeaKufabIILUj0AIHQt+87u7w7hwhXxymdvRAnuArhdbsB0N
Fa2cuOfBtmTsfQG+4vfpPajqU3XMCnSX8VlABbJkgPa5Dbm6G9H7bCERiRmDfg4cU+7G6TrtO2uy
bzBXIw1CUwBIv3OzIzFfjo7gJzd3BUgETteQuwOB8XoSu44KbYPv8Ni+cEI8aMvYzQmt3NA8WT/A
7YpRE0ytY3EF2ezDp7yLGp2qSNgH7L0zz0xE/HVk9iXpbJl5TpoAXKdAvujHG/mpqzk7hojoHNE9
uESFOt9gMVZdv2OtNUcunelexEH2w7pRuq/Ksrr0SPV1RLtJfDtvrEkD2TYguP5AnS9Bsb3ZMzMI
Wp8MDAkjr0eh4sApkLnnCuh1Mj1oe8LFnLt7OfZZGbeKskJZwIWs/IuEkMq1ga8X9Hxn7GkaFppg
liBj5zBQwbS3O9cdjbZFZLCsTsc00nLRkRe2cmuM7RhnqAkN9zovLBY7RTGFRQRMWM+PZ+7Kpx3z
7Yt3+LTo5rATHxAY9AzNPBJ3lm+Vm9l4HwnfW630t/V+cR7HBpCSWRn2o4vzBIy5ZeiB3yLvUdRQ
HSoHB/ciia+CP8NovAikVpwqgCS/4NUsA7NTsFrxB32kI6wij4ApJDSR9pCzRjrjPdx2U6H7f2Gi
fUnGPyKrUmf71DAxiELWzmZ6ehrpB05BS+4NYz7cxJ6ShNUbqPOIGjXitqG0t9TdmS9748hZaYM1
8UVEBMHZcM+yxPg4ReZOBpI+ZX6pW8eWCE4Go9kyrL1frb4wH/kdt+ftA+XHR7dNhQJAKOkm3eAb
43YNkVCgF92B5tqwd8AbOWclHknVOdv3NjCGJ0PDXFm2Wj/iuaReNIw+rSZzBmcYt5v9qAhIwf9H
EzzWRZdr8bfC7dYVz3cKSEqid+npa+kptIAMG2wqXYKPabwVWOJWHf1WlEpEqCBX3N2NpPZ4iAzy
571VsHEHhFECnmVq4wCwtHtOeAq6HV19I0jUQiYDAjIsyb1MCFuKuWYmm2Q0zFKnohHA8m4CPFK0
1fxFQEk+vYFVhXr9idUQhYXoYq3X77bkCsHv2d0bRhQ8y7EZL9UZ1NZp2DjH1YMVa9fbS7LzdKy7
R8MSWj1DqT7DK9AkNeafdAmuqpwRwM5jIPuX6qGhXVyfohqSGeTMZk1HYDvrGxzi+wTobXKPVmeK
bAx0b9CzHXbQJFXf3M4cC0wJbJcjjxgXKG9WFI3X+MyEDK5ec05f2nXL2lvIMeXoGarN4bAt3QPr
gnjH/Nqy6lpDGOoiG6KYJCzT+BHW05dFP29nC7z5aGrMknbZuS65jMyXIVrI2NxXMELBgDbbA27M
Qnd37MKjeDlbDf5B0sz2NRZG+HMA/NNwg7aRKwreJLhzdd11zaye8RsAtcMXYY3ZJQ2J7ok1VxwB
loZWJIleG5PplpJf9TMcN08V3L/6BS341zpADKEh7USjDQlqXnA8OGxlkNd/zHv6Tp10Bfp1n9C4
B+cJO6WQJ7gMPR6GL4aXSGMU6sfVEu5I+w1iai9g/Bi/Tqt2m6rADG3cmygqwxQbV+MDLKDNz0AS
sybrUCOXYJodHuil8POYDEEFpejr9x1nodUeg5qlQQx49wDivNXn7TOQcda7Aqk7Y26YBT15HFAi
Cdt78lBDfXU21uzJvExIOAkxJOHmiZXnkVT8F7Kvw1rUXcN07BJFv96pinaeH8MGilWjCn8+9oiT
FZ3a5m3x2ZNvHKOtBb3bOXf+tzi9Irx7Jclf2NdY54e2S7OP8F45iupCVrTEW4cK64vYLqbCPFnd
aR1BsUZjhlmDJHo/N5xL8nVRm1HyEnyBYvJVMUW9ijFcuGBkmAwqfPMeM4M0MjIDIn5Xe3phpx27
XmoO/C4IsXaRRvG/l8cM8ihcsE5tdL1G1E7iwnvTEOxlvdFOyAPgwcUDrtcObFElqgv4AaeEoZIB
dpcGq7nYYx7VN5oIWYJCxHj64yaTwm7HHaxsvTsG+Ax24MSk7vmyQbGaCCrBK/Pqvpw3VNH992XC
nGpBHZQnoJWYLRGBxopXtZpFYLcIKRgKJV+Pa9bZBcDgkZQyuVqpm4v6W/WZPKCpVhmGJsIcaee5
NAq3B3OYnK3cS69FClNpdsNm6PKfdPlBcm7BOQrr7kNzGB/ZPCoLdFnnJST5yGyHYPoy+w5bUuY1
b5B9+zRgjakq9Z17srldebNJdBWn76SJUN1YXiVxHzAxDA7vha9j0yYAEB1oPBwoCbn6F8A4WtBi
4Ahp9yIXBERYs7bOGVkc4S6HfUUM9TezKKAaKBKuCvUKFPo9QtLplTA8tbt29NZHXt8KbgXp/nuE
PIXXxjMgH9V/DAmcqrooPcSsp3+YbnoY21xP8QUZNli8e229IPJn4UGwiHb3CTzdpukIMG+nVKLj
+Mgyj4VraUNlCm4s1uG1+PAuKctRr4DkdsIG89siA+ziPFKbmzZ3EQGpqpmo7LKEGf5I/Gv1h0c8
hR6/0wfIggikDi3yo6Y/lFFIA8vnuxxCMyaYPCbMP3J/nnc79EKkBrl3BO2QLkeREBCPJH3RjTgo
yRLLLRjJknq5DsY4vPlaOp7fz/pIXN+ztd949DHp5BezA5eFgq3BXwRKTAx52tsCT0EiU2I0Xnqg
GssPvad7u+QeE9LPlh/UVG94uAessIBt3KN0miOTlU0BWAdO5kLb8iS1xFGuVv4hoBdzvqvKww9f
4B8b82K1FUgKO5xWuOqeTj2BdMyS8HY010tj5dN4sFuteAgoEvwN9CrIiXuUNVl370Rahr950Zbh
j3nVVhmRUR3K3gl62kfO0uHnVnbpYJTJtrwmNWvlN6PX/0VzM0yrsZoiufXEIzTaPkcu7wCr/xqO
VA+exRTZ/S65T+mgvNm5xnCWmNRpeGbPpmJ3GwoI8wx4ZOT47ltPKhWPC/ZNB429RtGTii3X76GK
XfOEndF+zxd6YbA5gT5FeEMqmJX/fZISvdqm8yVMtfZn1e10/ikXqievRZJVZIxD6zbMNRvgtnIg
rMX0LY0f+6QTpDgNvPmGNvEzY1hSkY7uvMPwHDhwFjXke9X6lah0QNLhg9Yn0RDXWh2hMjj4+mdl
a/OcFwzdPVEC2Ix9eT363Iomlr3KY013uVg/HTymcwLoXKCg//ppPupNolD97YrS/R2EEAeEEt29
XjU/SyXROnVu+iZmOrlZQKNGpPY51SirZ+NHookLgu1SspeVBzziXOYSstQLCCQ26OQQZu10aAFT
vjIgKagTAHrN+D+SK7UNagS/8MydSleLZb7XnpwS1wACjrFYKEk9IkDMFxo/Z4Tft6OY5JP+rYhu
d/hlqqwvXQr7WTpNptV/UzXzjlszDCIE6KnwBekXQnnRHohAVUCyoocmfA7lIWMv0QG4AK3457Cv
3bQJ7pfaWQmWV04A7cPtVezI7RdjLyI1sE1aOd45MH2v0DPQTuylC3jzo4fA2Aip1LUty7qrWtO8
dxIroB0ZkVriay1L86O/T7KGee3x+SZN6tjmuAKQTGVvH85fBm+i6ciWLFetmcI1xsJDXQuWdCvU
8w/SEhDZ+z0d1Cq6i3SAKb4rK5sGR243gwH0+G6E7ursbALRPqvwjUAP9hbKA6pcWHZGbbqVc5hC
lCY9W31kIMso4S/jRuENytaCjmpfgbsus55h71jalK+kKwkudp5E3er4t3Kc4JDrDcsoW4vsON3C
28NekjMAdVVwIDqJtPcCE9sSxYvlPbV+QjFuwJvoktL63gkCzz1o0y1ws/9zRyT7a+m6A+FMroVx
6fLft7W2yxHqDXRieUk047XDVCudizEhqPnwXbQbtuA8EVlPjD+k+oSCygiCor2UXN4ly1Hx6ogz
Urmlg7cFBH/6DxcUfDB8GclGiJrxVQG8wbX9yr3+E92RW4+cvcjdN6MjP6iaqmxUWjKaNRZVevKg
EkX6mB4Bn3rmKdJTmVHoJxbmPbd89R6D8CxAqyTjzfdTmQO/xQIRfn3RBXSczlIXKMpKpq4nyaux
p6nzcotJblwcQsMs/A1F9zjaKOjLVuvFpYnbVeiBd2M24rGUj8AbExcyqGV0ddkGs+BNLTN1aBku
/hS21znBEaIPlTsYBNOoxjHf5O+pduwkk0wH0piAiKp5q/Zat08x+bDN5zbO7CG5QU+/0wmNSg+Y
UrZightnke9vrEJ/3wuX9Rqrg70bc4CY5HlOg4/UvKm7sixsVjxdN6xledRDux/mww83SSaNwB8q
nLKnemC54alHsuh85LDFbSTqwpR2wGNtC3oZ45Bu5UCpfkpseYDTaC0AiArgJuyoN/jiFGnC31qH
Qbg6C/RYDXuGMXmr3NNii7H9Dhko4THtWCIMuXGlQh+tVgxEgAwD9G8DKXalCb5b4VtfibHV/Z80
JgV2P9sHXSiZH3Svx96nsfMBHRY8em+xO/skivPjnthnAEpPydgquAWQOY1Oa3TS4bAg+dZ/60vT
XvYLF7mKStQ29TTQf/uZ6F8ALY7kKhKEAmyoHtuqFpqv79+VJcmZyKQF6tKkqC4qTsmcxnWESee6
czp+8q5YhY4ZdFPGWJ4Mh4BMPaXl4Ih/q7N9or7sfNSdbui6ckpH7f0hciOB+DJI+czsiaim6c9+
ADkrIbFfQIra+X5WHHyabSGnsK93Wn4nGRyMx0KlZ9QKZOXtGosdH/FyYf4gxyaJp/WVZgCLwTBT
A/pM6a1NBBdRX9lfzUXnNo1p/xFJaRFoNQGPHtex2cCS0eUiQS9Rxj3YT+iR9AJLUzuqDhZl8pIW
GSA1Gr+ZoY29ygMWhgwCqJ7CIqMfjivpJsbaNavd4jGrH28YLI0S4TlnBMTgE2bvmtcewtdDj5Ie
26yV9yHVimPVBm+V9IS7HKzJ5DXIriz4JQCOKC1h+iE8cgx6ysaclsyBUD5EReMYhJtK62aXAXiU
Gyi5wzTExj2esm8MkaOpyLQdcn5ELA2fcKKCeiUY5okSD0JKLvKFuHEf9ZMNYXj/omGdgXJHFRN7
ZnNACbUqLWdp+IZZ7RY7HtTJrRTBus8IpOx8wpn6UHeTP95kKrH6XEpc3hk0LVh4xQB5g0XO66Oc
BV7FfPevkMIAErGewZxcg+YrAefi4IQV895f4R3h8N7EYqHX9R5UNpordI6SmrZaGd/4emlP9D0V
G1wf6LbtJudTdvOPAXcoYzbm8C+U7ER3Ob5++wL2dKAtdU5rs8mXpEEytex7sRyTHrZ2FNALkw90
3eo0hp0MpQ7dOGYSok8ZbRJ6DLeNyikv4YW8cXg98QHhAoaa6jw2r4kgykXs9RPMocToZeHMuhDc
RHdxY7kgLeMOyzcqjGSBxsp6KFUNi6QyWbWhtsZwk+YOQHfCLeONSJLWtEvoFFAGzwvgbeGM1ydq
IOfUO5cHkjmlhDc7K8wUU5lJ2q4pk6fQ9Cp1NTVgImCiPkr1xfp3DsHZ0gLWKEo+peP/oe43L1ti
WnViV893LuADtwHsdlcJeuR030UV+O8QOkqfdHtR8bJKWS8WNyVcI9OQyUDG0F8+Wy1/HfPLjaa3
CHoEl45P6ThM01oaYFM6pItsyiLbAeUXcrbI/vn8qE6pImIddJq0zSeO/HWyug/FvcNI7i9rO/4Y
+PDgQKxpeZfhUw0lFZZBG105qMHuXUb6IjP3xrcXpVkWnJ/F7BnLbVxHO9mdTT06Iln94xPkL/Vs
0ABA9bsJG/n1j3ETYXZgyOLFhKCr8nC9Qj8q8345cANbukQ9+z3AHOGdGWOEEdYV0cvV+MSoO5qU
1ff3xv8xdkWx9J6fvjyqJ8IHjFI51PutA/xmH0ysy/TqudTgryp1zj4DFmH8ihbNw6qc8Buzog4+
heg2Bz8zJHIxolKw6eOonRU2kjwgyuV9DWnCWJOLJVQHLKm4uuakmNtULd/PWPigdrgFS4/pjg1X
1CeXjWKNm5TmAiRoxmZhnIUzdIcXL9u1EjV5BTswvpNhxMg7GU4O8nKcEeetexj6jloQOOKkgh4m
5Jht+ncuWQ2pRc9rJ/IgEIgKLtvAHKsWAywUKJSnSiQLIaWYDVwTyLHacr7DPtWz7WVqJleppx4b
8wrHbgm9D9pYA93pVEwWNjxR9vOAGRrt5ftaX/PHtWl3qoD5LCtKxT7PD9qKJEIy6kfj16r7jp1G
PWxdVn1FNVqzC+QsBlXziRk4w+PtzyTzxhBnH0pKVoIUbbOmm/vxy8WA+oFMfxyo2k1atfXhQb/F
ew7xp/do6f7svIQRh8mri2uSIwwrPRtYuAPWhXALykyNH1hVW6ldcwGu6v2E4B+Ii5sDn3yBltFH
X8H0FodJINrWpJ7ylT+61W5/Em8WGE/dFd2XijJZL9cgMD1RfTPaQxKWyp2R2CmR1sm2JEmOZuq7
c7mUccpchiqtusRhhLUWfD3LGOxwvx8fyJ4vfZ6sxy1hg1iAEObxu2cT3NTtNKrX/kTMZkPgBqAJ
x61qYU05XeJynciqMDGJRbJoF+mOS1/UKt5lDFPL9anUUtp7LmdnUOh09uDLUQtgnJHCxtFnkHec
GJd850YVmqw/dTgDyvnnDqrmfMSM/9709+x2cRTcOCKuuriEeobc+aKICNROtV/xI1TCJzjxbyqq
JD9klFjEzs1zijTHBjh4cYkORxAwKltZEtImc7pDzVfzfrYagjtOqVUnPYxJIfXIGcEmyjJfQ9CI
DuR0Mks2qE1BZpCFrbbfkv39BPh6lbrpCo9PYICUtcBG2Xof4Vtgzp59Y0oa2dD/8ySIIVZNvoUa
YhvW8kmbG9Ve3qBrRprQ1sj4qjyBXJkL4O2+oViaWKMfTIA5eL1WHW/A3yCkqbGOzk7TYickIM0p
xmpX/iaFDwPSq9rUeqdQCLFQNobgDVTAKh3qkYWcbVpfYcGMXq1nxqsyx/J5LHl2qsSrmymS2W2o
RN/ZRwYN2uWcNKSK/TtaQzyVugXqYY5ckXP0su0K1rxqqwXXvz5xCmFgnvqo4BkXGDKieBu+kBA3
oZgkJTN/hb2t24Vc2Y3eZLD28tG3c0nGCFTyNVL8ylgOLet4uBiW24yVMMg1UHeFXppZAjitl6JT
Uoj8TgjTolOk3FuWT8irUpmR/uuczwXEeKQsHV9JbxLqVgUUKIsaH+V8dcyQXPpiIPlhD46tAFnh
+HcnPbC0fRgX+FEBOBL6bVS0eTKa67Uugj7/N8ZF1GpD2juP6RYOYeYEAqU5AuqqzgVkFOaRMW1M
m1kq4BJQUcZqxdlIebtSH5cL1ip1UmqVgAo0zKGpA020W308dQSO9dMHHOisBb0y6i0efEqZjZDI
GSmZ/d70ZChAQYGu7Z/8LQFP+z6X6PPSP4ylAGQWrxGl9rpKRgD+gA7AS7nz1ric0UFvdemNr1LN
aJoa0Ovg8UPW/dk0+oo4T+m4fgyOfLNtsTxB2ad0TPCGwH/s8OZT5PILErKVI6ghC4yFB/xUjTpE
6nM+TQQ4ewOjbAHn6WUKpevnOXPuB2YwJpFAfn3bC+Fib9hPF7zmxY22Zx/scioVzCPyJDcN3BHE
Q9hVBzY8kOwAthVUcY7N+mGYFsS3EsbIY4Xj88X6pnLjSQTvMC5QBnuuGbLFg3K7dmQzWopjA4Or
w4MRcvdxZMVd5thLLAH8tHRus1QNl01vKneOVtmSM8Dve/7HR6MBPvW6RwbEbc98SV5D8ZFdesZ6
UThl8fkRTH5RdGvxbkH1YhAwB6tbXIvzG+bXnUsHLkaETaa4OVo8MJcEQ8pWdGnUbXwRSwfGJw97
QFLV08ahTZpfLfEIMBq0GQheD+YH6+08JcPdONa7LTR35sVlF8st72D694yAXXY4Zd19cR0N88qq
r64iZknq7ZS706O7Uao867SwFZGZ4rpJJNKh0YSMHz65bN4WAisH7acDtMwJIAUiL27LrS8C1O9Z
988z/TDZ6KvzSBLp3Wn7EqAZFty1j+bv0Dopxdi6a/dS5sLJ9OnE9tMDMuDguseu9YVe/vmUQOkw
SBrh2kIS+hLxcwIYd26HYOxAFREoIuyL2x0XyWoMju1lVyNL8D2wKp5rhXZsSMFQZBJGLCeNdgD7
CrnEgmeGVLCBbGja9wOWwEJOWU+v20h1iML3JK5LCHhNx5uNQJQdj33hdsQxvpTXU2srBSaL9qz5
xF57kbQ1hSaA94aTr0jFztp63yQ5cryA565BXvd7RQEYDLPHTQK3Zy7Kxh7IsXgKlsiLUlAQJDER
i2uM8/UIlPX9gq7nVpTasdIipNj1iP8lI9U0XHY4MQXMp2AC2q8DuoONCcAL3hd1uj1CXjvrneTY
F2hTVrUhNxEelAFsxikfNaTUPt1i6pVRAjuKzxJ57u5GN74h96xOUipoTXPDPNFBpNhGuCuDSzh2
ZNDUk7y1vklBTtp1fk8fNWlvLz4/uB8Mveqs1PmvrcI6zHB4pjMcWHPWNHWNdf5eaDc1NqZHBqQY
37d4C6tl1RpNg3Ve4+k6EvltZa6P74DFD//pYfF/Z4w8XqNo+h3j9GxgoGA0OJmC1nKW62IwXRZz
w/U6PSm0faYeDbJwL197UEWtvl0lyIKcvgfpu9IR8WLEbv+1guXyfI1IappqTn0niXFQNKJKRGha
qnb9FDP2uC0Zuh74G5NggaLfC99psO9rIPyAPRFECilxWDrpdVXlmUBEZQXG74QDgeSjN5AdAOpe
+pHjSEFRPg8ei0mh/DtRGY3yneSQqtDvkO4rpifNzOJmRM1CZzKD9dQzqUmlve4p/pjOe1r0Y0v0
p9f25Yin1vrr05iEHikRDUS+j58PtQDZDJfSqRDFXx7vgHPWY8Bp6ZQtYtvzf+X00m0pjWR7Uk/4
2zLLSjfIUSm1qTh4wOxTqylTH6j012dwNHjNMH7g/UoCJgk3KPDYFFd3uFOuv5slZ/Ojeg09vbL9
xVQIK2WK23Dy8yT5qpsM0vtOH2calLMGF8Gqxlyia6o9TOTmFfio7ipO8K572UNII3uIKasXarC0
9gKmFN1At9EMbYg/GeOX9yRL2aCayCuuCfUriTRVX80GKcsYDJpnl54SVsMqct6VOWR4l/D1xTBl
sa2kaurNT7XPR024ePiH6SxzpP5jmvkLSJHZdvdbbRlgZddaQtbmwLojJMBHI7gchRtemyAq30DT
PXxJog+hUbRekkYGUy1thkZH9Nkt2qbxUhIkM52HeCUtLehJZ/TjEtoj6N7wHXOhxHg468yJ5NOL
9ga3Ftj+oreV6zvoQybpQrFYbI8r0ngycgDV9D3t28roNF+0uCuBQwQf7iO58ZFyyQgvK4JrFIzM
GIe3bduB1mVcKFmfO9LLpIQK0Q5Eut4df+C+TNMgKZHXp9TV/UQUS1IL5bRLB519g1hIpT53abSC
6vF3vPov1TdbeAm3TPu5xGCKM/ABJeW8aoRLa3lL/ujZKmHJ+y+us8svsF+Dst8WzO9RjnpNFOVZ
dGbV6JFUp0jgUqe15aqiv42IqXQZtv9+YpfIfxQAuBkWtp7PEXG4QkAJ7512Uf+rd50wwUPJ8ptH
Z7PIj8ym1Ft4n74RRcrNUzXdEzXOrvXQ7Mumm7yOheK2PqKkufBcvnPY+8+gnFSTed7w7ceW6147
+mgQzb6FkFepTWYyNfmG2K33bfZESZNvflptr2DMloNLWMaLq+3QpDWEUy5k7cMCoobLEfo/0BYx
i4WsV1kSGvMutDXTgM87/6Kp4U9NR1Z5HZ1eRQqTtlBPc/rMoCUlV4SqydfebAT0a3R6NRLGeOfA
QIyZxg5RJGznRlkuIxmVDfcnaT9Ceyl5muN9y9p5doqmKgx6tOq+/5LlpVd4OIOZAba6rvO4jswS
yh23BOnaRuvH97LVznN5PVulTMzDkx+qZW11Jb12OHkBMvfQ8YmVg13J36XZDQ5zeuz4Kfw3d+bS
fboG0hFoz1vlO7B1UqnlGFxugjX7iC2YCoIjDacTvPZjMQywM5gqt2JWbhDz/PurBMZRak74FPy/
FGSuiImi51UP6uFPIX9uSR3XQ0U+cf4DLP8aKmG7jRrQS7GKWGc9JDHOUGq7Ln259vOn1y8utlp3
Au4CirGETAXcCXDz7/FnzEYJUe226+Ob9p94SFxM7Iif/Jo1nlZ0CpDnCvGp5/plmcvA7kRkHOJ3
CEH+uvpmfWt2QLiPKEO569qRyqr0PDCWoQdk+pn8qVDxsXv9aIxzrfAA7r1cEE+KSt/FEsRq52dR
VVPDF1z8PzJwfmVcmOtrTLfh+adXp4GkqoaPWby8O6OAA0gnjKrMMVurdkgcsUAmlPehPtktCOBX
sn8voz6KQib0fu8pRcUdz/AB3Bou+g4TPYM4oksH94aKQTU5ACBJGzbBG23OzreQsjOPWZUfueEz
3bXw4KqpNx1P6LPN0QYqLTn0myhvcVcspVMdpqodE2ewQK8v0c+9CRd+PmwJI6xzQu1mdkvUkKAh
GkhDtLYKdisOuv0iYUAxYFdbFfkWCoxhG2fw+X6G4dJQyYuKEHUY6ko8ZeebsogE6jg+g5pVMIZe
IkkD5aq5qDqxmZ6eCytTn51SNa8Ivh5H/JwXpx7EqyyweG+LNu1dVjJaoa5qdaeeKCEp2Puoeghm
NFyHBUhkh9RWP1OtrGOyDGoO5Z6yOS+rCnkKJVTRnhEB/wAdcI/9s7WTAG3AuabWX/YWiuf1QES2
sfFeQ42z3X5f8j7XTvFwRGFAPY8yHoXpM51CdfralgrW4tHCUDwAhVvRWd8+aH0cUPiMYLjblzjC
WJjSOta2kttviWH0jXjdEp9yH6q9Mj5uGOWUvgNnpuAIk6OKRnlbGpJaVPyap9Qq9CjKGXqyDeeO
slGO2u4p2cpVgdMLN2V4yiPO2sWdtlHCJzikhFPRc+dGI+nyHjmASSkjPrLDckgQignDmEKIIJkr
3xo+ftbNUqz7Y8INx+98/AC686NQOGUpxuJwremTLV/n1qKwyiU3lbasqzpHmqFlY1OVjH7vZu70
y2sHQQqXKhEzMEgiXl3dswc7dIAccl613z/aDgnttGXZqWmpRpBtMrXcGLJrEEYDrHQBtoBzCJ+S
EyY1WIpey4Y9X3neP9IEORJ8IRffOrfB5iKtm7uR/Z+aBGPXwWruZgfqNMicU4/YA+3JGHvB8j9U
Pc9nM9kw+pKnOYGb05Bu/x/v1ogr+nCNglm6wHx89Me9oesTu7xhQfA8Y7p9G265uwP3PSmAIjqo
6T6FNUhMH+2KqwMRQu3avEiDEV1FctD8g8vezsd6tk2KXYZG6XNxCXrHquZBUaTbJbKWHjHksLLw
CB/Xc4hl1unBqhagicDy/71tQxujyK3RY/kAesz2gMIAGXkoiM3xwhNuR7q1njzdHrU/FFIFHnlS
LtrrhJc4BULDe7tY64HQzyQqECDErl4fWB5esevKuXaqrw1V3SMPs1wQSRrxBF4XpT3dMwILaWX9
Hqs4tOkmqTKWSf98HHh5CSa7nuKEDzQQNgMR6aFPv9yuNpqy0vC1QBiWZ8YGut+CZsiPesequ7uS
cvIfBVBaNiRdg1qf6zozbxGyf1/IFb7rTb7GVfsd6VQhkUSit1UuIMFOgUOUfjhI40BI8y0dsYwx
ZQtV9OWkTCs5VSFuJAFN+ffqFiDAXxMSWYVnX8Xacp/XIGLOaW2D06M4QfTlyIHf2F9Ia1ClGMep
0kKG+pERfyoKxeG78HFof+3OhITX4zL5PZTOcQviDIXGaK5M7YNQqG+ra8j1WHG4vOf66EavMlxp
CLzSJgLqxHACko2iE3Te0ykwrxgVzNc4QaQlTkE0DEfcWJoBt7Q9tbjX5hwSTVH+gmPYSfKEY7VQ
DPbw3DQ9JOiRC4rTnh3Q3DFoxV/f+4h5FRxg+tSIFOAbEgdMvlGrFFUjsPtMZCCvK4t/WgtkDW5M
i9fTXTO0MnYvpsEuiU32jqH1uahZKAUbbyDvmgcpII6kx2wLvuSVKiA17uuLRxIvBDAt2gPwm3pl
2geJ2cc719RzVAFrH9GbyPyjZ8saZ5jFoCFliqzzNTDtpdIj2LlE1dvAQuf1hpbMQ7Sk4fi+ITta
CBxHRXZ5Ne5yfJEpS6MMdDY070fjmcJV0BxBCfiLOLUgaazp5+L/r1mbclsJT3WNxjbvSPPAPH1e
r+FtXsZaaVzZpbyt5cvOqfSxJj7aLnCOSmlgiBaCxWOR/kXdIVPl+SVBeAaBuxj5EsC1b4//U6NF
oKXN24t/Vk0gFGnwJeqdjPpX20zQ0FxWSgt7liK+RpGKs+U3dbvu3I/infPZuyGr2mD1Ul2llYhz
Huhf8YEsaDx44kly0CQPi3729FxateUPHPCsN5DVn8iZmV49MUuTf2/19HE4yaqFSiHtFFXrghEY
pbrTE867ha3MhKAOREosfnfwT/nLNc/fDoq1dFvtRdIlQHjAp4t3R2jNbWS/+1/dmM5yj662cDt0
aCWbpBu6F/HSjQZCld8OseZ7VQTp7EjnwXIg26tLAvJ5GEKR9ZjL0JWY9kbXnJACrX9Bz/39Umde
/MYwwltSrdc//U4Wc6Kx1HRlodkaG9SHSvbOHN2+j7MrOsJBq5ee1pR0gkKVH1a3zTQYR/xCTken
Wg3FmAvwX0IUFbhBjOZMdzcWC4gDI/gS2Qq20atLR/DE3XyEdfHG5an9S4mY3wcFJE67GSYpatfb
wS6WnEAiA4rlollJp1P1jJuIqhumT22UjS69AW5gOC1bIHoqzrYUyyVIC84zMuTxUr4guuSyxhu1
1ganWbuXE112NDljOtPRgGDxx84DV3Tm4hLEjs6H4YQgEovv9PWHzIJ6OVPIT1ql2B2bd+JTGBLc
wz2jeKQIRotSNlEb1KfPWuqmhuSKdBll1ZDp+MAi9aIpi+lS6xEahitL2xTBhjIeQzU66PM06zwr
fEVqeHEmsmgd+ofrD/ugy5nodKgoYeJNGI9eIyvV+/KUFVEKqoU+DBZAHvdjNGbqqMcfXyPT0TUq
eCtGoYLvAn9Un1vhlKEGtmO0F0uj7iPqkjBOHZjHMHI92LhXz5P8FEJ/nALAbzci5Ax/E47pUmXZ
2g5IhRQA2zWu217I6j2X18Bh93TkP+Blcjm3mAtimcxQChYQOm3ibV3Ln0XZglscEB3ayfj+Qo+Z
yqI4odZFwzCRxBPKHiDPczUnDcJFJ4zuytbSVst4/h0EBQmzEoMHIHaeGpKQ+cCm2T3epr7wr74J
g2zFY6hiWAe9PLuMII3XvlR8l0JmG6fSBYQPLD0IviIRnOXcvueIftKCoIOnN4f1j0cT8qx/5Pph
vHSMMmKNNsAQWFVlM8n674SMn0xpYrrl8TAsoCXVxzIRK9oQUssJsgnMg3XWLOlTQJZWW3wQthXq
tGZLQLQ5VGbMyc/qF83b42/Qd0iOjGOd5l3kGUz/TU1wxLCAQRIQpFsUT5j0Xg09TBaD3NrET5Ck
C+K2UYUALRt/2BpCe8jY73sD1YR4fTj4I2HxVFMxAmPAPONXdQzVI3f24KDYxuMSj0nxd1igA1zK
JqBLvXsWBqC8wKGQcCUMMVarOjEDk+tJihbrOLxGH1TKZk+PmXr6eVq3aBVk1lJMz7twmGxO0RtK
5CnSL3mOUsNp2e9AWkAPkgXCqIlZ31M5IwucAQ3G/Z9kHRhcspcoIx0Wjj8mnrzkdeOI2YnUr4NR
wrNJLHdiuqbkp/owACFA3crarCVx/0RaCKA5c1rnBnnQGFjyzktG1ABkHqRA9esGyF1aNfPTHNsV
g8jxAA6yc/CwoWfg81mx4swg+15WNPf2XuhnE1G+0qaxfH9FAQZ6XOnw2xbyuL4cKfrd0M3uAhbQ
XugNc/4KmsJAwh13KSlc7C6rwU5oGeBKocQaOPsLHEW8YLl9CRJdnTrAriBTnp7SpPQfw/o4s5f6
fX0m40R0I+0xtrS62u6JUCrGbTET9B9MelaBtep7V66IiGBUhzpF+9ZEntsEKnEUldvRzctPYo21
xvTSGOrnMlVSlU9wvEdnwVyEP6M7V/ft/oeMtMhamn93X/Fp4sY5XdALDA9a2Q84WJsKW+XicslS
cU1VL10xqaf0sI/Vtj4/OxB64h26qxRrMP6NDGdczW4aHIrTj7FbDRT0NmS+Ve5ZWlM3aYjBS6CA
jdi70YjtNZjuRkEDEKzB1MLTjycGSuEk3p3yBKMlhhZFJ5D6i9rnJACwb4AE8WAUlgaMyYdijtHW
MCmdfMYhq/EdUIBlxronymBKBoRINJ/KB1tuHw/zFslKsIuUQGwSOtrlq1cr91RpafEuEuSlVtxv
rXyYKbCCp1y2l4+x2EZdABSORWEMM3TohMdT9adGCYHnYOfTIcFDa8LZTis39aVQPZWvdfJbEukc
Cji3DW+QvH+Bj4E1tXTy83rq6jQ9Lt++fiS8d4GGWPxyEIRHfQD/IbGEU1HKkbLo6JQOG6ZijdZf
+O/zyqzd12RuZny13pldY96M6hbHp6TKMkLPUlHJRkMVbHEyBCCIUc8Gy4ILoKPkBmXBCku4ihSW
AXPSiIWUA272UAjac3iSHBAkxgafJblf3ddgxbieC/6NmxmdTx7tXhF5nc7kVzmxNmkT/PFLP6Zh
H8GLE43OJeUQXyQZaUSL4UZAYWDJDziMVE0IaiBI4YS4KD7nwIHguhLpXgUgSeDG31Wwphf8A0Ex
t2mcHurXbQfavpHSe8JfpaY2CsvjGBq3VT0j+48hxGQwKPE3Ov0WbLgQUtiCCxyPH9+vLKacuD9T
pg0c1pwf9jC1kVqupuETpwstJtxZ/hxeYnKo35NblFCZtnjtkjfEHOAzmYTkHTooWhGFzPP0HcWH
2KJQEi4reC3jq1wCyA5ogEOd1LPUzxXD9DTm2eqggmgcgX7/fkfU6+zjIvaEy4N/TjJ2jjm9l3YH
s4sLLZLklll81TvmQ02++an/746+AYv0ThXwUK57Z/CA1eWPRZaAn862kAJnV0ERLT+ZCNhBMJtC
T9eRE0GZgtnV6mPSVvY9menfBUv7EJo8rzL84Be93nfiEDB5kTfpnQceps966yibiKkI/txSMeWT
rs7CYpfF1rR/JQ7Yu8BLfxV1tVlhgBobNuRrQeJVk9PhZqwhdFfU93DrR/K7U1dxsrelQLvO6J8i
drd7K4c4KtT/TEuF/qbOfsIlWGvaDnPAuZVGObTQitQ+u4nnjrQ9Gv3oK7ZYezxrY3mfiuclk9Ax
sVfQybB8B1mY2Y1BJqhNgecAjPC2XXitRcHkxE974vgDP3D0Yjaw/iEPcdg/iBRkTlv/0ZJHv5+s
EgwlwtJA49sO328RoCkn7wQVNg3C5FuWFvVZhQCctoZ2AKiQnJrgqnkZKQp5RNetqXcAEg+ageRN
aZCIEsJrVtZSaPTv21zu/KNbq7h81tM8xqu6T+X6CzQg7UUZmBB3zFveRs+CrVZdj/dNREkwZYnz
J2pbNi595jxNP143CinzXQOQDpMXjUtLcDiWYgMkev6WI3MmYN/MMcPj5vYCszIixqCvP1SWlb9L
4cRrPa2vDk+ksWgqMjRDh+1BDGA9DCSFyp/UDgMOEyKZVt12Vmho6jUf9A2c3Nw/DtQcbSEmwEKL
OLjag6tx4hx7cTgzxrqJ3vz7Us68Pxe4f81mAgo8zsYuKYD1d7KOl2lZDV5mfFHXS6fR0hihLP2l
SlR8TiTpVOk8wVz/SNZGbTjPLSOzW3SJi/Vxlqg7Oh2vc3yEHCGI5Vpn2FOiilOF93g0XG8wHRQT
HL6ClJs9/9oJV2OgJso2tVcjTOgSt9s4iUi0byHTnsklR0dcQLTiYt+5f4zvQnMZFsOmUbHnmV/a
Wb2f7MyI8Ii47VojjNphhRLgj6VBBnDoYOBJe7FJA/M/Od1e+qn7/ei3urm4ylWX6XE0oqMUQlMg
qs9QxI9UP/NWNARf+T9+ES/DfmT3TWZD5jIV8M1522tmbGgCup9XrKbrPvUkFx5/43NdfuA3RAkI
R9Qfg6xv3k6IhefNoDQAFKHgavwss8fV2fsZtXzZoEkb0yGhtrT56v2K4AN2PCGLwzsiEp9ixjWD
7eKSxhbBpxmA+HPIUisRsBIH1/lDefu2J8IE50wORLWX/L9iJC4Kym511XgHD12T0+bp9Kj+AFHF
kLtXYsnfkBupKsc2SpoC1+9+6mJxEKtDgU/urft0X3wUe4k5IsTIJ5tNx791HJLZ34xlsXOSMnrq
rtyuLoeUDlM1LnacJ5it4tT336FwVJ0s9LGjiMn5tQJU501Y2oNm0kinG3vmXiu4T/5XYNttXoxW
9lrejzKtDurzG0XUPUuylEDsYurGblTq4owyuMMgnH/+kQtmP5wuywaWaQrs6PNQKc6+W17UJdLa
GCmYu7LJKXXu8GplFnxhYvz8IBJqwPgqSjg7pjPQwSeyCfMUxs+DpxDCG+blZCSwIZtlFTDq+jlJ
N2nUgq8BR3Gz8zZPvQ5xiUBI5XObZ9xXPoVSwb0AJzeRCLE0eZxE+aopuTW5Ys/bVkLi8aJ5CJbi
Ynf34m+t6bzX3muHInKJd6UAf+nww1eMicKXBr58BCNZtN9xiAx+tbzpIcwvXQmyrFGOE4fadthv
Jq07U28lArI2CU/caG2hD7mJxkD2I1G5x/eHEHaiOeOqKGCG1HGLT6Jk1h1krYiPnOfoLOW+g00F
HTrsIHzTVIwfEhTImD8yTyS/5WXmSWqUiEz/0WlWdGd8tTN0D+Yw9v1531//P1UeMrMtlphb5bdB
MjWZ49qMXQFdMVT2EGC+lEFDzCe3GxmdhoBe8w0Ccgh60H9BnlLx1uuyoGcx2Ua0cMvjdI8Gdhxf
MjIM4ZCCgK/cVs6QVCdmp+QuFplqmDCtVn7wb455F2vluW88nJR1BN3GFyGb8okFoSI8aeTV8gw8
cQo05ZvB3VWkPvbxXZIfXR3wuE700MNNZEO8nvmqWiENJKLjIxwHOdj1Cc4zr1jBFTZza5mRIiJC
Yr/Bbd08fAmZX8vpbEdjjEVaSSxTVokAkqLV2HeK7pCecYy/yxGoi7ROh9i1AkYiPGcMqzMPR8yv
YMKE8BDt+t8qTd4MbymkBlitoDzf2g+hbYA5EYSbGBfIDptdI31Bot7nyt0z/kyWvKJO9ufJ2EAQ
jkEmmo+r0uMPrpP/ezIAPYwt7CsudxDDG8AyqWMpA9CXCG2eBh+kGtiCkMZBtnXXQ2h2yMAB/0ms
cu5D64J3d6ynPVLL/JI2164A7X5I2RQRgL9WQfnng5sW/kVwnZ4Ghlw+Ur0dGJDLy4/+L+ITFYu7
gTsMMPT2QYtttgzvaQAAWD3iILlGPqwrasg8wTj0BU+UWCH34fU52ZGxboToH0ZB5MqbgSXnkihL
T/ya857r1MFMrvGNZ/JVLwzMLRX9PWvyIipOWDLPKMNKoq+8Zq07+185MvZXhwcPYRDKvPBr9zAd
dkrxlo9iMBBq2alNuiN/Syo72gwJDk5+dareSo3xyB2VtiDv34XbqoXKr4/xiyh1IoPlQytm/Gh7
ymWX1w4TqxPwRNrdqCEKD87RhUKOaIR56i2T9XuQBbosRqBpzt6P6/VV5FxiMirBB8GY4yJAckZF
U6RcU2X3kyFhegJaJ4Xn+/qSokprQLdvm1XLVnkFSvLwUS4yvFBZL7o4VbCXPIVCObOTrDZpQCZD
9ENoGLdRWky4Uxw12/QqzJkg686T09LDw2OQhk9wDecmcXYSzyI+LGgT3+3KPjspQX4VtDcY+oDE
o4mMDT1RA5a2Walk+ix6Y+N2V7zaCWB83E9ck1kQ/dC4AGRUewSHWZxTp3+XSrkZqk3B5MIYwwBX
oqNDKybj5Ej2GV2FF/d/3zOq0o4fb3eYAc8dsV3sk9DFytWn7dx3I6Cm9iXsnUYs0/hapt+YxvMM
DMZzRSAyibuwnSQ/Up2WPImJ34AvLDknPADv/P4kutLGz3x1ApSXhS71/j/sNDTtjp7lVy57Onxz
yNUqSsdMew/kEJHhEOo3+WSS3uPUrNB3qC7ytMm/13dM+1kUnmMikFrHL11xBsaIdZXtmv9w0rkR
4KSLE5elqGKYCNT46CBM1ia6b9rPANivuVKtxBbcYXKX+URs19tD4sU8BNPZYmWKSp1S2UZyeHZ9
nQmElDkWgA/dVhPhrpoEKqiiMuj6LrwGoKoiVMnBY0wRmy9JH8lxQetqjrEievahJttAf5rzUN1b
YT6Q0rJtx64femU1GOGBUxyDtKp8rmWCJ05CF6f0qut9LYKIVQyLjPI7RLrJgOcRR0uInVECZRqa
u38LFKi648s3Z8ShwdTdaPCpwvA7P0Pmgk9ezkgy64pJoBLS+jUD+LSICsh7HoP99YBK0UA9rsa8
nb/O8pc9RGwdiLF6Tjjkvx7/vKyerzEiSvgenPQGI3pNurX8rZxx259aqPNWmD+WceHVitmTjHKE
PxCOYNHSR+OUr1Jhu60Rtvim5DAzTnC8u+KZ7OONKrBHIk8Sp4+UpaoSiS/jhLbvLWbQFFRUqsc8
SQqrDiPe/Q82MYNd4vjktY3NaVOVx6DXzb7eupZmiLxAAfzZUzvO1HZtSZXrqhlPOlMle5s15+DU
DCRm9Aqa/QqM3oCD9TXqSINSRfgzkQ3SCR0/Y/h47Eo4AMffp6jbMb/gd/0qc0pJvMaplkjVITIX
dESmINDVCX0rfUa7E7K228PvhuHdCUop2uTT9LrZNpzdEG0hmJKm3E+5hYIO02a0K195ASY6DeUK
CaD9hulcBu4SqEFRNjs2fN3IMNf1D3TuN8ugGgtFXZb8CQ2GG2iI+PXdQe2RkxgB8xcvt5Lf/Wpz
fxVRxLz6mo+AZpQ8lM/kwQlw9wfqjh8TuIpMXlbXdssg6QiPpK6S7peal9/hN5H8qzg0gBDO6Q2V
KQ7eCgAs62ByC7+Sa9c3fgg9b0DlsGI1jRBqLY+VyuqZK92yHveX/0fwreA6lg34W3OJez3tqKrH
9OZoNgFy2NF6iTbmyhH4tR7AZ79uBgPSsH2Fs2YDsEWt7v9If0xb270CJHiDsTpXx61SwGyd2Ldv
HEeEzSrnS+KnD00U23cWMZeek3VVc7uHtLkRgPcsVAkPRH1KET8WHL6Ch6xY0rmKA3qlSDRZ+5U9
mitBC8vAoTJ/X89XUCMcfPdr5Qc1vNsyLxmmEkPiMNzCsjRrFx9fcgVrC4t5xkwGr1zSmqh737oT
5EpS4JpVgdJ9X9q/ySqTsafbYPrRk0fWHFAHxkklrtzSnslY3z7bnTntgpp6r5xhwvk29bjpedgz
1gfGfR2zQZtMjK0e8x0adf4bKh2EDemKkSflOaEUxGH0/T2UTHUDxh9BbPzaeDAlVZnBgxLhTp3Z
AroYQNIuFlMHlZ6Q+53xejexxVEQP0Vcc8EkthOGFxRotSpS+SB+F8bcExh8/tcXluYTn6TZNcN3
s5nJiEQhLJH6jS9ud9dW2mRQvvGcDXdu8Y1WKeFLMJdZUgUTeB/9OOXb5Knxrz3DZRJsNWEvVCaa
6bV3IhENbkkFDfq0+/CI2eSDNN3caNEPyz0KYMne6sZl17KuVHFcmJNTCIPdTlHmdcGZjk8C2Gl5
Gt2GRIYzj2OJzwpccyK86xvjQ1ui1AfbyIUzoPlk5TwDJ0Uu7P/6TS0atLJk9gYcGxwIhauMWYWn
mdEHEoZSDapkNxkx+36kE5j2XvQChAqs4f3E822AfgQkZb/jS1cw0yOBAc97fIv4w7Z6ptCzPfJT
C9X88pYC15R+htLR8il7hw4DMgkjKHusmUghFZM9w7W+RWsYzDcBettWELouHNa/8RzFbgXP+KKX
bXqVTxtBsXUdssiHOLowCGTY1LSZABHV86xAZO6hI/dy/W5T+8aOgu9KdorSEHJnpOXQRkvk3M21
JxOwSQk2HZIdLghQvF5jX9tfqXa+IQJpenGqZ1tBlXhd1HEem6AKYxUAsNs5ORFZuQH4Ccgek6Yi
bHlaHJwMylZG/19N3ayKiqQoSqtgWG3HaapAONuBe0EtRVnTqeHQHxTnoK6U4uGDdwCzI6XMlilO
2R4nrMdj7oLFSgHf1ZwlV+swTPXXLh0yI4+U/cjjkCI5zw6iDLkScjRrEWW61gH/aJF17/M8aIyG
o3PcaPR33rkpBb6CGYQhkgDLcr4pQzaMuHD4TptigncKi8LmhoJtOrIQWSFcU34OlkOoWpGHmnOy
fz7qoFK2H+mvV2mOYNBcqUDE4IgcPbOy0eUcMlGN7cdVTIN6Li6WhBJ9gPLteEaul4mHGnEcRJsv
kQ4WnkSxOuLqnJm9VJmKc7W2RxNsmbaBbBq35GlMDPG8ljVwD/3XocfFFdpf6yEpfimCuoPgEThf
AtWIUhkKAtPx7VI8i0rXjghjTFCkzOfgEPN/qcVyguPyZ9US6pVd4VOinLiY37j7Qgw5VjIl0SS9
nmSOGyzUvONIvJq+yEJrZo1nSWbBGmJLjzI54UwmTxWA46+KBjjC898QzLxt8Uz4JbJUjonKCYtJ
i/EM9M33DlzF7Dewb2bnQrKDQsUohTiaQlXhXajmDoxseA+bl2dTS4vyYCDI3sjN93y8wfdJy/eE
nj4M4+oxIIYjR5/OOgzO5F/8p3SHdvwmEEX1cqWkGn7mN1uxuwuE25l9q31lS3aU3oS7dUtWfrYh
0HykK/u1DIHjDQXfzFWhre4fhgkjcE9FMCV38NMZ6OZcnEWcNz/oi/n6Az0swkOPR4zXCA1fDNaE
lUbtCJZ5tgK4k4Ljk2FjNz4SZkDi/WiX/955vQT08l/q978S5EoLsL7JKXAMP9Da9b8TP7gkuuPs
nlK9XHbYFozCvvBr+MUNaoLs7D0SZyltV+IfVrxsBTZrzXa91zcY6Rfr1FhTXQk7pC5Y5EZS50KF
EwDgBv/jsQnDTn1z8EVMdFIclNniuMLwjVlwzidnjGVDG9wwBukmN1RVzVRHtmVgH3A5A6TmKXc9
omExg8JJBUV8iI+RKkJ5r6rbErFV/TMPGVu99h1vw3YmntRhtutFnINP++C3Qdz5QxWz8U+Qx/a6
QBoTwBK9HNp5um2/qp/NZd1H4UdQVrjtgziIfxskR4TEhtAHI4q3SvcS/Z0/uXFnToM+fSxt1och
B+WQEJ7uLa2khEh9ZsFGBLc1ewSUbK3clxOPqIP5STKFa6U0LkRRdS69N9d6j9B+jE2Vzt8oRb5z
y5TO7V2w75yfLzdnb4l+JYbDtzXHnPLMToAc36LOc29x1EdkDiqqJ0XPgIUpm5GPV8AmfKJ4snbL
MSn36w9UOn7bDLAjfktKKqGyYos8b14G+CiR4AWppc+9pIDySpUztTYk4YQ3TWk3s2WTdS4drQs/
51SR8f7EDmrb/q5uSQsMFo9LMISSDH2GcJeTi+vq7BV5bjgTA1mr7sGiqeGdos67iHQryTx2tf7g
JatDDJXjPdukHEAE98XlcNgUCrPSJwoWC9uDtyKFgCuts6pBaCeNfwcvjYtswO6qJ2CFMpNc48rr
2+lp+HyD34mpughyx1n4JciDKrWX4J6ykkH70/sNRIQjR1+8zXGQXDvQuh+wE61j/B+Qgc1NHQ0B
BXU9EKAGWedBQlZbtjTTimXHwfnRgLqA4DoUwdnbqXEQVTbZtIsG9H6pPzJrlmURTBE7MH71Y58t
jOzPKlet45sTxrvYQtHiEVpZyB0ScGOZ5TkrAm+ZPCufzlrDWJO9zqgxSe3pQH+x8sG1Lgn3VSVy
qdORLo7MSILtPfL4gHESCoV996D4Zx0OaQ5qdkAryc6SnHWuRHy4ozkpjoSwI2JfqtQ4fCDlzNsE
qCiJY+Edt4lf5N3fmvx9YiIJBhJNXhAlY9FRtkb58UVbv8Olx4GhXoRZ5zCD5Ob2NBe+FqWqjnoy
G89wBdLefEsnFMUFjWVIFSc2oAhmkKHyCRH5WM/q1Qy5Ji2GQ6az57wJ4AJ7zrrIVaWrAM6+YXjR
GTv4iGUdx/it7JIXld9BilH7xoM4MToCut79hGb13I3WncfiAjrOrd03HdBwRqueld1xJIIvrerP
FvEmbE19X4MoVJY3c5RQRINAezyTiBJbUA6UeizTiocrwkjqXWZqy3/UikWH3U6V1eaEZU27OJau
lRyRXAoB61JMBvcyCfZ+NwfqKTlLDRjffh32LetBbgc9EklQiCuoUA==
`protect end_protected
