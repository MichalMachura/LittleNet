`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VAgno8OxoF4iBvt805EvZ5B04t7vIuHc5hRCNc4uRUsaMd36oBh//VCaV+glO4HOAC6/d4L7akyM
NoqkXUiS6w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U6ZhtQdIHr1gLfhADEiO+K1WNlHhBgQb8eYI5f5jFHZ5UYXiHVsQATY/FbHqztSmNPvp4KvUkhej
thDIDPlHNW8wgk6+SiKuMewlbnM0hTFcqlQxhzGKVGJnjKT8FZJSPSGw2Hg7E6qEHzgbrJGQTlKF
73SCv5eKc0S9XMUe+YI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NmFaPLOI1NIvYWxm2v2L84T3lWokDxeL3knkGbSe5KXlTRb6J5Y74MKblG5cGKXhtxEkCQ0gec5D
hqLTIc3UcPyDzE1CXLtOuKOsBoDPLXY9MKGjOCgHy7Go+8BDylOwPYNRiHe/vnCxO7wyHu57IT1n
pgKFaw/pAxxzchjSmQe1RPSco53iMrHLJejXCc2nHeGQn83fPc2bpT0Cq3aLpd12nTZ48EO9v6kO
i9G72xIcuCkS2V2nXFQ+dv6r92AFFTNsfyQYpa6sHmH/qiOtYlUIFoPC9HJOjFONJBkrwAxng/DR
3jHngCh+/ffUm+7Y9cujnFzZ/aTAnoVqDkUJLw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tY1Yr8H3ZMvW9KPKsXgsB+/u+HwJaMnptw8PQcv01FdZa0ncpM2nnHZPwinabKiMlgHSon8rYa+C
BuljUFY8uS79ceRHr5tppm/0ZSAiSeWwP7WlAAIsHzXc/f7eSvvJWSLvsu+zT2eNJQf+wFqQyxJV
TngIxT6zxk4Bwd0va4YF1lLQSXA7fpgtiOihGZfZynIzKvD9VR6ua30wMSEJypDxGdHtMD+A32e7
nqR4FuqLBuvVK1JyatqAcxGXOVp1A2fHajEnqf5NCIT2o4QU+h6smFJ4pwfz6yReEitw7rUksNPi
DrMGoh01+VaYBqSmUHllQ9D8o+qu44747/shHg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
epgfLpE4AfaebCd/xo6rzntRHWndFcvWv7NNzkC0DrGgLx/qLMeiAzPXT1KZrOlkKYar4Oev0KS2
seAzBZKOJb+dfLMfGjbNjZPeLrLums2ERTJ7WE+5yAv4QGFHxcC1k80l0qUDCLHzBzVXW0c8sX+B
LHmVbu2gMQx5y1FOKug=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HcfaoEBWp1R0frrTjXqZyqFBlPGNyaVQrS04wcexFhFLzPM8UsUlXJRxmZojF+CsQtP9tf3acyOK
p5jS6LsVRYWE4J7kOtXgjf2nKzQ/pzre30c7X8lSwCbmxWMlSP1GufuOv5x4dSTTbF1qb9ZRy8UQ
LbVBev7PH63xB4SwUZtwkVYAh7W3p/loLE25DWiS2Qq+ppB+u3VtZcoVjGoW5dDbqJ8FsAJDXNx9
hK0iOW8J5gFbMT4etSZeXmzjY0pEI7idEQb0lyKow5bU9tNclcqoPqqopsi2kqNhMsVaCpxOJOdD
sbnpMAwKMFjh7exSwv5qauPaTMgxp+RfABM9jw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WB4hP6JlC0o0M8+Od+R3rCSDwZOlSfXOLohbHV5nesvh55O8sjA7b7ir3feizh1nRYijfKi8zTA/
WyECFs6xWiRGtvpNafeKuhORfQusbndgqqN8HDpwLXcpkqymf4ftNAKIgzUlHIPOJ8Mi+NzI3N8A
rjYnA6wkoBCjJn9MxGPgJISSjAVsoKFBvb4Aa4SV68hp9QqLWlIrtNajJq2yl0w9O1PlvObfPjHI
N02/wUmym0wqIfKBfl1lCKLd8yZRoWw0AwV3EMX7NMr8VDVwpp1zuxEMXX5zg1L41p1yrxXhARAG
DgsFDrr6Z1iW3LJ8ES/gxOinFkqrootk9Y+8iA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VN0xOp0nWW+D5ex5VOj6GzvPAsqIRZ4LgrZZGNGpxBfhf4pq9cO0Ptn4shsfC1tVOJ9LkHwp+FsV
4eFMXd7kWb4Y5GG8tMrKRo8Wj6MScYwE3JsRvi/r0c70rq05H/iwvDN6FRkAk25vpinAdfiMNHmp
KaguMbyP+OWVsWvL73uCOy8tFg8SjkQe/MKWOROFyMOr7+5zxCQK+pDmacX1Pm7lKNVegyLD01K0
UeYpLhDeRMANFVPv+dHCtKkh7stihgtk9qfNK9NAFg/JTmDcfvs2rBywQ+S8svu7MNBFUuwHy8AU
w4Tor65k368a75R2ewdiua6MNJgvTXqQ/XpM8A==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KX0I33YSxvGDPd/LhoPFxFV0GNRAII5wmVcxqYL+WLsG+br/lj8z8lthZeJ9h9uPYthgpfC9Ttam
D/b0yECdgRL02fw5ZI5v9XZTb3RsAMXY5DlfTGsywmtHIerFQLVM9HR4qDOjVL1ATRPpN9pgNDbY
HRpOKe1JhvtZWGm8abiIqzYoxkhVZdsqld88SkD+EgjC6QXhObic6fdS1A3J8xaLHlzhNua9/fRp
1pyw6iHAfizbz3L8vmEwfh4uCSJ8kmuDirAAZjDm7U0OjWtp2MYP5koly1f526/KdtukdtfEkJVU
N7c02FLMvcFZz8EzZURZJ2XCKAElKtQzIC0pbA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 271984)
`protect data_block
U6USm8MyaG9ScQxrsVlXFloh1sKBbBJvFvs9wIdws/W4R39KQp9nk1HjfExPuBFbVUWSoDWUKSKi
BiGfyC7I5KwHobQgFCTg+d/rdAlH02qCZfTeOEeTeqGT714VU8TcCGDUy8Kmvk9kFE2SpnTRUFPo
NE8eTtWbI3kYZzWz7LXfkWmacWVS8cg7FxxJz5q53C3Cdqs8cJv23fPDJRNgxexrzhjd8/kKO5Ow
mseVWIM2/IwGpgc/o8Nqj8bYRfUCyTMMh3vdi8Nq8TgekLs7/ZMAS0PlhMhQo4TY5k2lDkGJnDCh
LLZ0Ah8KarHFSaGOINNMlZqd+YwfEDDBeGn1yK6JtVv9DW9p8f0pNr8ilymY8FlBoa2dRT+FSYew
GuZIqDRrphgfygaGsTvJQxyVuFReZ7XmfOkF1Kj+f187wZhKdSn5Mdxrr0bNTgQmTG4RkyPXdTtL
suTh1KQNTUBP/p8sApXzneiSOO6GxWDw2jxFSLbHHV5LOspEE1CUn4htlMiYxhnyVdyLbGFsnWzf
+O+W489GTvhtuGt0npyXxwUsmBTQuPaiXJDRrGsp4nI2BZRD2+DmPuIK/5jsH0V1u1MDOOBxvgAF
sWRvlstyp7uwtNTDLrfJqD7v+t+zTgLoec5Rd7eLmwEKeWBKyq+/PY4s/hAj/l9H4gncQbxruqGC
jRMNezjYFPZGeIIELZCZ6hDlvjIi8sq9gZcsDsgAfKPBeOAwdtZ8uH870qblF9tLcY7Qym/iZ9+M
leNCyvgpZ23XX5MtLOGy3St9UlSweKycHTf/xBORhuF7z7tibvD/KcnVqFJ89bdTkmbthGWxSNwg
KRuBEuQhQNnLxjPAePTX8rl5at6jTUfliRJq+5HSk1MjfcySY5uB9SEZsunZGMKZHxaBhZrWtG5l
d83od8WZs6XCO1om/GYyZ095jx+FdSZ54FPSo8qjvcsAyHEcemf3GE7ChoUujXoFdZOjdjtGW5e2
IfrfQ8n8LnXix7YKopydiW3zP/k5gCw0pc5deLzEoNMc4tBDoXMIighCIjTr1nWbkJcv4iAaATOy
Yt+GuidQRehRjW9ZqhUeNCUX65sp4uHY+zv4fEOxVo9TBjtQ0MjJp2yMn8ptNZBbPsw6az844HOY
7ACW+SqHW6poJoCiFzqbMY4pERzJ8H+BflhcIlsuYEaPzhKvYY3uoGfTF31p7/XrSH2VGuivw/tL
bbgAYa3OeAnZrIwB8N442OEUwOb7g9YsNLEnbs+qIqS7u6Qq6B/OghjZUQ52nD/g2lciElkmLzRh
wszfN63ZgZcmOv4YxEkRcbRTSBPmNrDyn1M7DDa14HJjQdkcD6RZt6Bh7xorGBWp6StUNZHwqc/+
7V7FK1+7ihV62h5ZbZ9G6eF/+zMjzpydTnKzsBmaJdo70faVSVZLuQ3CK0wXsShRDgTVuGxdl6nQ
aHf8SY/ajkCzEBuSa22UYsvLRSELIEFjmVrDXnG2ikKEGK7I+fG76uuT3Tr7lIjuBkOPpEojClz+
UMdUETsWUU8fPfgWbkqAQuk5sMomVmkg/CH3pJQQ2Gxl9gHoiov1EqFKIInzsoqNlHbtsifjoB1K
vySir8Ksvz4YvpxV2PW2QlAb1ejkeMczi1yPzy+FWAhADYh5Oh/3JdnzuBJZ80rQMbqbLb4gGyxC
SLOa8dEWB7RRSXOZwYW3eCaa0k0qSLWe5Pv2DduV+1sZwtX4+NGUjIk0UZVvBnlp7B7hRpzY1YG8
qjnPIikxsDH53hZDARvTH+HxOspAsaPB3w1fkBSChsBuHpP25sOF4FWmFv4b/BSecahiSYt4dhUi
aYNhYf0aoXbGijyH59vebOy8z91pUPCKaKJt956n7TFRMJHQ4AjRb8Z/kujkLhsGaEc/NkNWuwvs
Qv5ZcaboeAhO6bdFipOsOZzc69Y1W+gKi4Au/Ip7JKd0CAkK5RJ0eplh4m2aqMEYLdABbFFyn9lv
XhLdAnWIS65pTiWB24/crqOBB5p7vMLqXzokP4Vkj9wH7HNbxG3Zv60UqMNDOD943OPVHYsxbTz0
WJ/PeuneG2Vr4cfVVB87H/Oi+ZwAN46WZGOJtRflhZUSF2jXjUsqNViqsMFMD80HXnrre5B7hCr2
fdGaFDt6vmGgRVVB9jVhYCyR2Cm1QsP+4SuhbqTdLPyODtDrBsL+PijWrAEGetrcDv4bkuqP8NSs
sptoG8fa+AqqjrI5a7DpoYKumBxpC3EF7Sdtk2QkC0FYjL0/Y/nJzKFxkjExgGsEhFkmov4YvdYM
WUzyv4qU00HE5fCHOwqzjsxcYuH+v9VWBOs5sp4xyenlrfl75G2/84XvbYap9slLx1tgk+S6x1UP
D8EnBPBtGPW8Ejs5qIbop+lPrEbGda+V3noXkT3j3vTIc9o+MyNLQiVfb8Lwa3dIcUIt/ITVhzuY
Yv/vHTKUuYv1MgTAYBpG6YwAtf3z+Glker1/FPDOVzuKFUxtUbYZEZVhmzg8isIWHl8ITdbDSKvU
adHNO69YrxwS/Sc6i3d1P6XvdbV4JiWB5fx4JOxrqVUmro6nYgGH1koxPoYuyd3RJ4H5BdZEkEv+
ZzFi9uuBaODYjxWq8k7b03JtSd5KThYS9wjH72dGuDS5ezITqpifl51w2JsxxWj6GLrRHX6yhBQc
fNbvon86Q2UCXNbPxEjdtDzspKS0z2su9sZjVs75zO1q1jj/ikOEI1Z0lH3OcYpsMEEzyGRN15wN
WWZedeieMH4oUxj1JbA9c3I0IvuqqQ3Kr1JcpkJf+EaS4+2Y/IIb0AyIlEugF08Rq++LGLZRuFjR
/xlstebF8wQbt7uBR6d3dPLHt3N7rcMJYs+UbDkxfxj+YGNAe4az6DyzLv9yXzdQjRSSaPZEk6qI
dHx9YmoDc+mM2SUZZsUBFzPjFOHIRlSCpWKKXx3Z4aDd/mQ9iEoDp+KkpN4yLct0QA/D6poBfu3F
yppymBPjo+2vjGmUPShRpgaqsCE4zSg2UvUaqJ/XpARXYXY6Vl/Iyt/CYhHJJzS3vQM5pa4KKDWk
rsQxsK26rcOFsMgHFz/JtO+XdeIcGvJXYig2KKExzCKVOZCodz0nQyiw0e+WODn223l3Rp5u5F+j
2WkzZWf/FaOY+Y+/awNdmdOzCyu2RnTyaMOiivFJmbRKG+OZ36Q192/ybfO4WP7PhaD/SZ+Q9TAz
kkF2A+CHIi1ZjexXf/6u88zbe7sGzY/oW75Uu2SgEla3YW9ew8qrvB5v2dxdrqn1LOTaEnImtP7l
bPdirx6YcB0z7ht1CjYw5EZqz2ye/5qvexq7JaR/zacv6QSLNP0b0XGTb8xgKSZ+XiHtWYjtjccq
6gclHskopfZtVmBE/NtMSMGLQQEttfc+WwZqpgipdv9fbqQmL16Brt/dO1TpHm3QMH+Uw/A3qV3D
98U/sZUl1XnuuatUQXbyWKIf85BWC+kfP1OrkAnmWDukDfoSuV+IuTa2MYZoaU3LVdzMuhYf4Z5b
b+eAT3lRy1dp23/4KTk+Him3/+gfn+3aSRhJ2VNkvAdPAQzq3IpQt0ec9voDJE+WRn/lQJZNsxp/
5EHRRz0FQRq7O8rsuamsjk3+lWZ5rbrKFCIAVoyBv40pAHWOGNCTQkdgWccuBqlBIwnz0U0nc1dV
iAGcphvodb23xh9SCgTsRQoUmMP8NHTD46MSTT/5CWd1JPxAoCPBShq1HWi36xM8WmjMnQtvh+6r
5lYSIX7qd8UTEoZCtzROkjMVCKHHitB1z6xKZn9mFHEE9iI3po921bpf2n+402ng0s9RF8vqNR/W
hWWalUipW6VTn/kFqNGSgVMKQp/1wr2v5xGQcDTZweoJ/cVBf8IhBY/aKbbGdWBworGhfJplJ7ta
T7KZexFkKFbWTWeqlP0nRTclbv73vVh2GmvqYZ1FtdiTCnhi9y+pNunyPlZ0qGhNRXOv9nwwPZgt
g4stW1nImNN2N4q6JG17r3qN4h+I5h0v4yCcqDrT6zJMCx60jOVPMoN4kt1R6Jvy/Qb8OrMIpfV4
cqGv4eLWHEh/gCzKqzHk9SBrDEVNoTZ/mXZoFM1K4H2dfvq8d7vJh4sJMxTfJs9zFSYvSUQW4WTL
wEJMs5d0Zaw/tqrREc0MxFFLeGLmK0BUZ4mD5ua9kWZJsz1kzo9OoI51+L7wIBo7Gyu/hQpRRTKr
FbRsAyHyprZuq8eBkepT8s/KVI6Hpu6o7NuRkZU98IElUX13lc3udFJ9rZP1JvMo/F/cfLsWVR4r
uHPCdEzlI6rwE3Vghd5WMSQ8dfmsFajQCplzI+xlv0JEynrKOa2FNCkJQXmnTazt6gg+8TxQmTxN
1+ntVz+EL/SMzVondn9tc/zk9EEGoj2nOw3RvV2atqPGuRF4TKJcE/womCYog6In83vxyge265gI
B/7Ca4SMCSBiw8pogAKpQ5+jf74n2aYa961oBhafxOAWxplESHUZmo0efYx0shH215BI1XY1dwfO
st8riXNg8AQYzgb3YRsbLixxE23sFhtgHONRlLopvVJmsQNsF7boe4T3GznK+Bc/b4Rz/laGKpP2
Rue4zKxt33LWt/7IIWb/QSZ6SK39kV8jzwh1YN8ZCkaHL3ras4eRZyBNQRWUo1A5yfQDjlXiAzJ+
agwmw8UWucvl/XF/60lTz7dYxPRGX44PlQYZ9swN4li4mamffY2wmSyziLcoiJmuwSPJOVNgPCq1
mxKqNKbgweFARVnir5DKF6ex3izSdCGaHzqEsLuiEH+uG0OA/YXWu9lJRd0CFE54o3SvvCapRhZm
GG7qufOQFd4/G5niytdDG7brsD5hEqAexCVAYRe2N02X4NlJApMbNlRoQNoKzBkcHAQYtybma/mH
o3djZrXXzlL9TnxTlTAWKQQ3XOlbfH0QQKxvRY+AkIqbELOt7ze0VaxQHBw02Y0G2cMrtKRryQnB
NiSPDjQ117lqAdfwGNWMuahoLoNb6IQHYbfD+0TA7V5MVnCSF7W/W5Kjy39wi0cfqUS5/YRppEiC
Kh0z2mL36aDmQ3hwqVialUH+pdogaUEAct/tYv+7mBhQcndoTjDWQoanE+5ZiEDbz4IwyxIEyKyv
SrYnzJLEso6hioYv7WVWANBDYWP5T4JII0yDkQ26+df2Sd2H8HnRqUrckWgLbP6/2maHxft3tyIV
7eplnadfy3NiwtCwMPO/oS1F4dI5rfRIZW87mDkSvUwq6vyk+WYXLmhrOaIM7uuFshMFapSfPmc2
dLDpGBspcHQ0yRbfO8ogKKBH2aogWz7uJ/qxmCEhPGlNxQ92YBpCu3AEw387I2X2NMPfFFNZIPlM
MuAjeSyh3sN3O47uUxOcfACMy20XCEfuXMHq5WsRrYUAg2Bi+XWGAsHgTCD7FLPhE5wjn9MvuyFC
A27RbtwO35NiWCQvhgzCWlco6cD8fxAVb3cv3zJT9Jp2xHL1oHThfgUvr1s1lAEjDl8nHspb0SZF
KY/5X4vahWU7vNZM4klw/pIGqiSl83Ho5NcYBznF9MdnT9XqqFXH6IoxwqIJcg2nLb097P0oQiOo
nrTWBCUNaatutlHYKSgtzjDRNE7sSPquaIaMRew7u2rulZgC8ddowFmgWZ1GoihryzwTpGGBtJQV
ZGzelMKmuDUYXNAmnlm0lEOyQj0tsYFk1KxeLyI3fTuaeX1apLmGVq1dVmPEOwDJfyhx+F+6V806
QH5HL9LUxBDtpZLutfgbZWcmukSVvCxzhxFQ2KW8SDmXGJGCeniuuXH1f7/FCRTzp2smiLMUciIR
B4+BpRJRnqRFRC/Hz+pAMf2SG4Wv+uDmCMViOTJ4JRbIJb2g2Oa1q214SomFgBo/Yd1qoJxHPAFn
8bCiUX2aQEfLBad9ieRC8h9gEbCDHQm87/0hdTeuaNGjNcD10SJPOCB7iwleFnkO70wRudVuOwhp
bdkJ+rBM8uX5Gjy0u4GWe9DWlUc74XR2csUNyZ8gAx4/jr1MROvraCTCT70WlSznQg2t0QJcVm3Z
e7TehG0ZHwC9VK6RcW3iccro0uTLpGe1U1LsYjRtOWwEVwUUh88yJfyFy6+zEwFHWJ9fFfLDQd40
PTceeUOT6vEF05Q6sfzMbIUIvMSDekx9BisvP3fpmyvsK8/xR+cW35pDo3fz/Hh6trYs6unw0pQ/
KNh5Q1T5wy0SeiBRIWt41aqTg/zne0VnG+J2F3KNZLWbABYnP6BiQwIKDCvJ67l+i9tlLV9bzB0E
cIGIpSFSUNcaAa1rid0y1qFVMXKXvBEzL6d3NhPf478aiCZ5Ra4H0lMRsOe+2hXNhTql0edqn887
vS+48ybKoGTm8emzjamiphh/1GfMoPlWO62plhTjX6S6v8isOabBCUnwLF3VDn7IF4VyYJkSGy34
0bQMXCzfw3Ja9ZJcRi7gWD2upRfBwHXKIjFmURNIJXaysTRoxgAtlj1HpSuFQ4c+khcIsE+fAdeI
X8jv/9RPjnLmMSFh8UoZQ9NyRTgR/BxqA9E34DKzNS8VHprZedhTd5mX5Io73TLSNBreamswQT2X
PnDPI+1JV32Mqf4lrcPadlJ02AA6z/04iSDHseKAJ1//53lm+ABnOnI2Z9R6IAhrHfKwi96YwTi9
whSwS56X655NVmfyuG2xtPPmGpdH/6O8piBZTersvbcOmQYqKylJuzdNxbT+B/OzB7WgzXrgV3iK
9JhvMKtOOlJaBMAbeQ+lp27KlnRScXvdLBCM01RRzgQnILVR5ooaFlLUDGIc17mYZeecDlk6xYXW
yhi7TXv6PRF7pBmTa98yP1C9a79zF9mVaY50HuDnhxjE0pV3r/18HCnMpxZOdfkq6CbH3ntDYJYf
f7yyffADiWuTCBof+/3c6Ewev7+pW9FbTe58MPP4EQtn7Zrqv/tc+CXumiLRgh2ibGVopBqw2Xx/
soOKUQTg5lr+gMy5Qn+7dyo4PjKhXK8JBQ+zqyVnLK5XFGcjnoM7W4drjdvSP95VOxyjxJos/LPd
yBOkaXFuFRGSaM9fG2wOSDpdkuLin3DGkw+7EWKp+hIbFErl4L+lpuehFfJMhMFEm3atcaQIRo7r
Oc7BXq+nYp3LRG4Y/PGi0eW0s0f2uQNWxgAPgPNnIcTOY/nh9YAF75pYXSVg+Ijs2OmjLewhn+oo
OTlYRjeSYlahonXLpjDCFFuLppsmfVbDzQSUaeUjvxoqZ8IjpBNFyvQpTWUK3C+YBvyJjieMIbfe
WLompuEtGYYp3PAXdIILAyfC9uAO7argEj3uNX4UjCa7ZcPJNRnOpR5QtHvZ935lWRJi444UBum9
56rGxYUrJNPYB+EaCSLfaz9mah8xTQMTlHVcQOQmWkL0FsZcdjuvBRicnCnoeNVwoJfEwN4LVOiQ
vTaqS90Uz+ANAogaevH9jVLjPa5AA3t/f6gF0wyM8691wXiSwNiBAop8NdP7oJDfN8sgYBLK/aOO
GV4ZcQBq5uNKy21sb76tXyIvQIw6wYNCM5SdA3haIH81STor0dKFis8A82WNlM5kytItPabwVWIb
I29pKS+VH4Bmbi7GST0Dd8zD0Teiu5eZgRqUTdlISp9M/tBT4xDFNuV6Mnyv6LtdXVNj1HqCjhzx
RWTxIXSs+vR6G3KzGrQQqO0s5St+DpmLw6ztyiTkA7rY9w0zarj5V2z6GpC7a1bykJ2Iifw+B5qa
2S2dDX4yw6md+Kps1nvSDav9sNUEGTePsEWQUtHPE1jdw7dlTx0zqs/y7dLAGM0OYicu29UYN0yE
mcyyg2hnztn0sTTSKDyvtxp+/IIrraHxoL/Bi4KMw/BLV/mk+kmbTprHnOotO+y/a8yKPEwSHhaX
pEviGOB28cWpR19/0/ENRpYk2Rf5zQq8KNJKBcAnXCe0M9TCviJ7B8Dm8TccAukrXAG9DKjtapNL
YJ2JAMXU68/ULFBCliwkeZL6XqJj6QzTQUT9ioqHdX/4zqROyfiayy2qCPCOrNlWZuF4DyZO7jKF
A59n5ep1LYoyfHTKIaLIsTi/Sm3EfmxLkyU2j1MnbLzMftQuD8ffqjL9EmIeZXlaESjvXgVmkLFh
OYpQ8DHG2hUSecNharfwjUXP/lcbx9ppJCoqecZE3s74gg8RtLe2D+FnpZH6GS82lCePJt0Wcgry
Tj8IYSfGg6ysIjMkVqblqBZiEZvUyblZXS28+XjBmK+J/zJqouDjqI5c+6wZQKiU5crynsuoiWhn
YcaLb/dHqiQHSGV+rA62X5upXgppmiwXjP95GzKlkJ0JR1PUs/1Yl1rwymuFX9VmunKEMnXVXNZo
jMGsEJKqzk3SDh+wbWROAV2wBNkfK2e6WitRrVjAfQAg0j4p2jwQNCXtbVXE1HwfCpZdR/I6LOW3
6UuxI0lMihnELLbVfoG/5NavHUf5MYniyUmtslD2twPNyb9Lf4uxZ+vuSQ2Dx0TdAs2YxcqPrlK5
TW05B3HSCY/3Lv0ozhao+JkkI4Rf8sMuGh2wUWVaANhx/7Jv+eZ1iSjntAfP6EGItBg83/qT0JM6
8exPcYcOzNjVPVMwmoo31KfXd1kMD2trIWTs4F4p5gNzY+ITAXj4lVxITFZ7mBzK7FZ50r17oo8w
K6F1ffy+QDPEdE5DBK0fJ8lKHrFmmfZ5oLCvIO/4aVUmkXv2FXfxqiDgJEOJnAxnA0GUy1oc82Bw
GTUYmeOtTGBPUp7ZFLhYS904lVvB+Cf6XTWLtAHiF2t6WbQzbl+Hy0lCZ6DT+daF7Cyg6ZEkZv0w
Dcd4v/pnsbnOVWWrOm4tAxGhv1O9t0OwRZh75Wg8hhTtn0/g2gkT37OQ36T5fgsIA0zYztRZxw2g
S+VV/oIUsPWPzPQGeKp4RZhJSItD7jmMt+sueWZ6+943iJIVQorB9/xcM10F5YkuBm85kLKsMiMd
lmbv4Q0JhMzV7dW6+G2ZBhj0B7o3VqQWqjYT6BmJs8e3FGpu2bP9K3GwXkPl7O1olM6a0Q0HNu9/
/1yXl9nun+gBO1uc8IHPE6glD20vBAb64BUDgbh9dXFv5fow+qDrXTHfUTS1xU0gRmO0N9FVoSFs
5EfVabfcNnfBip/XBcFbFajSAbslxZ9Y1zICt6OUz9ehl24yW930awsu6GVOsWkMAvK7Rrc+W0PP
+m6Vg7IhixDgKH66VZlSN74P4sfR3I1FWx6BdjGgANhQCiwJ+bdHV1thF10WYvQ2UmHWiBhy5bdI
xPv+0yMwWfXgkgTX6+WAl6TyduD513oCqGvrd2GL5bKVYfLA1413UXOeDu9e9WXYwpciu5Vtg0hH
gdp8DhsWSxslNSAhv9IwhgTaqYv8cEQSw90CgtoNL/HN64h0H4pNyf6rSZ8LxYt/kMm7fJA8c002
ARcxlsvl4cSoT5Zb9k0489HNeDsZTE5S1L01H2qIDyW5Aa9lneSTt2D1ajh9z4dF6zHkHETN5+UN
0cc4gWsq3NOA/MZrb+QRVG74PcdxvODRkLyiyzVvhhpaC98rLVhi9wfUg9Lxls8DTU5HGrtYlP0o
wsIgxX9imCAkN/VnGMyZAh67xyVJFaUlgqiWeNAQpDAVZBgZSiLfGNjFliO462BOUNpD80SYTH4v
wgDJuX49QPt5ikG3NcIxYfdCC4oj4B72odkBhvtpXIqtsJU9cUqSMZ4DAtucURDhByrf59PO3hsu
gwMg18OxTixkqA8j8ym90euCw433NmstnK/jYPtoZFse7DSLqqbA3+DEt/mftAENHdEVsOJhDDRv
+xcYk4A5g1UjC34VPsUzPvRI847SEawMu0LtSXi5E5w17jdp58C6pm1QRwFwC0kivnD9Zo7C4y3I
hIqobRw4ATnkOcv3OBfFS0BxjaugRnK7G/g6PRhwmUh0Ufmh3hZ71HLYc0CPOP2YDtDRByQ0xHYE
H4K1EpmYIh1UUFVaY5v2ta7PFucKB+VNWWyuLQ3qCC2nqjQonIR2I+VirBOkJncZxVGnZARS/JqW
eRtl5FlGM34RWYXABo8VMIoMJpws7/kYoTMYFD+gF1yg7a+pSK8S6u1xQw0FWNMSsxoIrCQV6Bgs
nPX3LJ32XFmdKoSvu4PwVb7rsHvF9TzMIEmPD8XD0vs2/eZ4/w3aXaWEXpyNXwPyLFghtODFsdR4
PX4jlWVOkGXX5bj9GS25aK7jgoHCq+On6FocQANZNHvsOPqIFBnxAQZAR5rjFXlQUj4Trn66fZt7
9G74WjhOKDXBGrVt8lBfvq53GIRiY3VEzYvp4ZxoczrwC+qSd6L7zyiKNqCu6PDrgYTJjDT4mVK2
nAOhMsko6IsG+nMbpoJ66M/FwdOjPbJd5T8d89mz+hYEOy3QJXqHgvVqdwtOGJLnrPaw7WjERfus
dwJM5r6NbpY1kVI+m2RvKnGNNRxadGZDd+aYmzNU1BNvs7BnDUtI0SxBF2Sb7rmn9n2SFTtXqqIK
8vWDFBELJCtjfWJ1Mo/MhxIPoN0B0akpBHTmQSSkv+4hQczifIC6A08Xz0zQ0LwV8m8gjUmIP+2V
UDqwEpDoUyL7FQ7xvnre1xUBAy7uFOMl/WgIfmQKbRdr2854sG4e40qxIuv+6wk0LVEGUMm0Crdt
hG8BxaKCDGQl3Kb3VBMCBoxPxRAAA0hWEn48XYQeYK9EtkGyIu41nTmeuivd1cyfwwdqvZGCzJ2o
cupaW2fSg4KVyaeZQmRPKWy8+4Chtmi+xOpMEsUuoSsqKl0x8bGsF+VC9MphDLVwfsWYDTIdkgXZ
gGk2acM5OVEOY3LRjV+w2LOnfvWCzgoHZBOKV/6EeMPIgSmO+VpjrZIu0ElNxR/++SzoCorHeJXe
pgz5a7jwZCFYowEtCMqIdItPC97Ax7JTInVaUoIIrUxJSCoCw4nrSUomhA7k6v+cyxS1REKhBeQD
hioC4eHgUXJdLcp1LdXw5wReMBwmrgMRWYYkA4VNZZ9FEi1r0BM6khZYqA7ztA4wc57oKLT2iHEF
J6trJdT8HBEWRPjsOQVyInrZPB5aGG1SeP5/OjNnswGNwMzrf3M8FLhx/hfUgUZuDB6iFVTIx+qh
2GmyOz2IoMdn1XOI+wPB++VhkextK4/NpKW5R1KZFihjsqklse6QTyAj7sMpduckVqI+ZvPrABP5
8d4sF42sXDSihmK3Q1smFiswq9QUoNrnsKUA/O43l589D6U7hkgf8cxKrky+dy12H+HD5L2+KUB4
oRTYe4FS6KJ767RuwnTRgWsXUbK8IPo9KDsB/XAvPipdk0wYo3XOy5tELzufLQEQ1RgF8+G4l5zL
OCyL3+JbOXk7iTcC74L0Gs/LwbeAoKlPSTZOv+v7E/Y8oxUrY35xAKpOZprPFPt26hh9eD8+D90G
n0Y4FXL2KzDb9vWd+HzZIhDAeOUJ6+8YsLj6RJXI6g3U50jz2qOwNQ5M9kB7WM+r5z0rACVYbtOG
O9dQzfLZog/ikagoXsnvnpBV1kyW0Nu2Uuh1GBIHgSQmwRL7it3CXGJVgN5cCKfDC8uBO+unflXz
iJ49p7EBD9SqL+0/8dSfZSbugIftrClaSNUKD/57I2NMTgp125RQzhtM9MpGFglEVE4qeKmSsZzt
E/+E3tCmMJH7sP9Q8PS8qneQg3ft4TjZ6mH2kg0iNp6dXfQ93Kb5buEZF6mqAOwb+dmp5eT9FH4K
wl1u2qH5orAaD2nU/laKyajovRyPjgMsYiXJe4M8hgC8GhRJeaC6XlHQdkarFOoVYALhDCVo721n
/94LXTGl9UEecv+SVx0ZXh7URplmASF0x25UNufJl3O19/nUEG1XGoiG29fpqEW0LYiLRCIvy5Fp
xyX8G2m9LFeU/izbKGQN0n1/4jTJBlWzfa376QYvjO+YJZBsXmW0tVW9nRZLLyZ82eaWLzO/9Crh
MF0i9uqI5SPzd4LMuhrfFXk8xzDe3cSkZp+Cv/36pd+hXY5vqS5fE0nlL/tJsScfh/JhHGViwlev
dzrMELg5+fF5PkC/BP1CiVYpgCIms3rqtsllr1grvundc9lv/CmZqq9PSGB7yxhLnB8f5Z5ZwVl6
HVwBwfgEIZF5otv/f9TSxxLE2GwfMx90eBOyaKqlBhKD4y2PeivK8FA1cy6XXpaXyF9xLTaI7OS2
iXk8qxmXLeiRgeVKMaRD8/7huhiF+6ktQau2m/oei58CvcgMoGDJtAAr3xECiOAxz8iXW3tQ8Jbf
UnatwwbKn7T2uiV9Rt+xvYpR0g2S+qM+5ngw8o0a6MB8PIrNhu3yo9VfA8OAMbkd7pzwftL+Htm4
miztO7MPoQq4URE9u90zWJzAGVGiSMZitJrXRBq3dCnYp0Yin+gj0vDEFCUOnbMCzeqsIfrKWOV7
MDnMPLNqO6k9o3stObIC3ElXGhULNiK9VF/TM/h/+pmrD7C4frBW1RrrRCryylZ28KZkis2c21Li
EqHl+UkeDrMzszTtvB+Fgh6ggFXUAEc4XWZtPe4Vu0cwodnYegYGwcGaZyQRoBAI7M8otww/cnW/
bVDEoOmn5XdW185pJLBC5VBOKHU/WqQFY0OYj7VM8CkjBj5ETZsA8v/kVHJlWitctRkEZgiVUNhb
biTR5rAFcn6otqCXGHVRclkstDw86aZMXLKP4j+5S6VZ4Ff1zrnpZqIa6W6P3snwTtH3VnDeUQg7
ncoJpi2J55yYIzmkhMFvqJlIolNkQw1l7OL1BfvuIkPJN8hTCYnv7TdEhl50RQoC5lizKhZ+1QtL
y1bsH1W8vNKvKeOBFn3SJ0xEF1FK4eZtMtoJ5QXwHf9lIKYG5s9QzOB/P2TXEZ6fuA7uLvsWPrwM
uUQMsk7oDPS43yRAZYRiZUEPSLgCUoHc+C0hvPquIl1uOM4aUefvoENuhf/MfzVH7z3X4cssgjjX
7n6C8DxAdpkAPVHNaGHMuLqEQePhhBJxuzmOLZl+veCCu+cySyOlW09IZ+We8hXDqYCpXHd0zKuO
p07fhXXG4AYEbchbBz4FPD+gQe+YiKVOKhMB2Wy+gkmEaw+IkZgVOHdRtsGKm3gNck6HRfOBt9Lm
w549blV1RC34ztSLKjoGdg0x7EesoXSBEOlrM6YZsM3RBH6UEAN6brmc7WvWKVUnfyQ05Klo5Ntl
HEdTHFIZBvv3+glfvYsZCFF/1R/uaMkhavNUkNvl76DiREvrJmCM6OdAcKQYIDnIPSHmI/C8cUee
riCgdWFxag3Ndu+l51kOTrh8uV7GIjG4yNextzP4PtF/nw8A9u8aWLsR/E/W6feivaHclryKkoqv
OVpjAyqiHtbrl8Gf6ZrK6g0UEVdWGRDUhsdew/s7CiodbFZw8lazqXxWjqHx5xnmyCelptDBcLmv
Zf8wtqsHS220ijUPXH1Uolnmrl146tSC0b3nAVmMiciYmEJT8IjMzXHOB/TovxQ39YWsvzMR2uSQ
JdTus7lunamXW0WoSGs4Kj7DUVqkq4tZ8LB8iTEMapmp3vg7vERk4YW6W3avCUq30zBvm5zZgmHq
Lt0IadY1u/O+aS7Yig7THleEkiyfIAs55lSchcp/+kdnjtA+8PURe2Xbnl7GG1lNnIGMz6GWUQ8+
TQCfg98XYtfFP2jCicko2VEyaGOSJKxjrU4cuUO4piQm06thQQphByA3nZS0T/gDz8ByIQIenFdR
FlVirIARZ7T4HO+0GhcpWk+7OD/fBCePUUeujHsssPpx35mnAXBKajnI6BCbyltmvQjaSCiOo3/R
q8UFBuFKzZSb0jSNJ2T6jRPvDfIgC2dI8tR1DTNhcyHFW63FVmBMzRpx0/CkMsRKvzqh5UkGrXP7
eUmSpEAZ/z7S57zz0t3bhWjfAkLhE2h7WyGhsKOKz5lRl5wNXmmNyl3Wvn2xKbrAAJykTQe1yxa1
FrlM5JDLOM5Bw/FHcO1MSmxXQnDLsnBJXS37nthYBgbA7VaZNdbwRC5ERaiW4SL0S9bq8IoOysuO
CCEOTuso54z13tzVyfv19WkCOAwtrhcNzNfGQxd+X7ykR8+OjyAP4ksAk6YQAv9ZvA3VOfya/9hV
eFWyXc3GINVxkFMKSC02gnl0fwWNDHCyyjfzsdvLpjG/RiSEOUWb5bPBP9q/NfWa4btIXqwghw3u
BOWoiEVrvBghSTHi9Fp1JX5HG4piCNlhYib6BdtUwVPyx8Nv7WsqF01CL/HlCcnsssHETr3gRO5W
1fS41ts2mpp4rtWgfuHes2B/Q48neAm09wQ8EDdKDX57SXDxDLOKQeqppD0ONUiMsO/s8EZRLwnB
Z2U/CR8g0x6SV8bJNtpBVmmEM6RNj0qp3oCpjGHKqDtvz8UH0tn0vMbYpzeBg06CyAzF2Fny+eC8
GoOafcmhr3tZuhcjCyjP+J5smRdVuHDY01NLU9zD03wNMPQEQlI7X7aobiOcUPuzm+N3WD36xPON
rfhXUBEk6zXm0cDkcU1utyNSkkXOPBGLNcXnKujwzc2EKl9jZHuN57UJEBATo/lf1qczg7M2fdmy
7jBZcB6/Qve4DngZW+AqBgq76FWJXDb7r7sJdutSP5ffeRWuge0rMsHNn3b9P2GoU+vhaZ+REYA/
+ghBQY3/dyuBFsSeIS/QJCC19vnz2M7ObxvmdIko2vAJS/xKEhs6AAwNPkpOftnRwo/mRck1+G/Y
/Csk9e+XiT11SKqp5ZP4XomfjlUpb8ItnLoMWeleUPRyXY+fyj5XKw+/r4O3FbiS1jKITkXMV2EB
5iBkBzFt4uldXsXts7BfGkgarAOG8zhlFjeyitcaxfEFbjRqIdQ1+Y+3VGOKoEtiTdmDT6cFCbt8
dXGXjA1TH2CZlx0cY80khj04F1HwfMkGEDwaxjWul7V0TCf/iSrhvewjb21w5mpTk43Gn/4o+qUp
MDEBg5XwsBIWNFUvqMfGrKwK5A3oBljCiMnyCwfGAoLQMWhy4aAfXYuz09OepBB9wAlUju9AzYcO
WJ65QvwZGFlA29ahoTZDoGNzwkfHsvU4lATf15PHpbBOGaR+2yYCg1uDTTqg27QSanKxqr7TYVG9
eleGzAvUCguejU1yNJW12sJhnZ5wIAeMsXZJ5mE19sxi2bRId/YGkie+ZY8E1BoNo7Ez89C50fft
UNDCwEq2Ufb2PAFaq/CwhCOfj/xAIfxy/NxPI7ymWMuWs1hfveKHmzl8cr7WvO4gc1duS9jIl1Fu
tusmKYgPpr3haZVf/tvhRuqLhY+YzB1rhelU7xErC6rldwdyM/VqrNXqYFyIf0zj5ZJ26ty0VZMl
y9/tIJSv3oMZ3kU5hvFyUBBoMj+Ue/8QDbMXa5teFI/M8sNFpH9Sr3CiK+SAscn6SuutViHcl3qk
iv6uJqODPo0dqJX2FnuX8qRMpgcR4+u8ar52qYwBwQEDed6t2VeV9xjpB05/9OJfFzQwVPTuj/U4
l8Dk8uATAw460VvdwX1jLf81V/JOS52xpQ/P9qrItTHqLO30mODhO4yeTurrj3vYUgC8WKiGx4rF
2r63+qNuJJCGUBHkHrjW/V+evWzhu74F1GyJqsH5y/l603A2e9gi5OqIUIMDCPBODU/XiI14p9aQ
40puoEpDyF7sKHZCGLJd+GjrDCf/WaDdAkMxaVRSkhSnSktn2uoiV8AYkzHb8P0HbvhMDdshALVn
0+b/Ir0ShFuujia+FH74yGPFrvJgCKpweLcA+PHC9eG+9nsPI4NQO2d5RVtkCtMnSYEX9F2CsBFs
otCXMshFGIswXjd5xFJVkEjtgDiBeoHKodbrtQCxBPdFE66neMprFBH3xsAhkI43gdtW7wpZIl71
Kb3UKG0uxtJs4DnuelJ0KW3dHxftmCwYoq6htSc6Lo3t/6n0kFoCFDUcIEjQfbS2J7sBt+eNYOwa
qe/sGieP5aD/fcTB6it1rCJLTX/8J3yk51TqmYgFFG2Guc3BDnWR5VWDvl3a5HQ/ppjY3RGVYc+d
2zBubdj1E5KURDphNTz1C5ZTVMFJvppjuuPxQheerlfOnODPHPPlhOnQueXuGvRUf6uWVPjIfOQI
OAK2fZJ2cHPwsHKJj7mVL2yw3uByhAw7mFW+JOoas8rpmFiTlUSKw9oJ4F0aTWKzXJ5C42nRTsc7
e0vGnLq8pFZwqXIjtmmloxc2IrLvguogaqHuh3WmOloZPZIzDEP+GRVhFaGUHrTr8L+A+Ze0rBtm
GfvC1EY9gWv9vSWeQDMmVHj0b7ensktB7Tkhy0PyIJs9QYyLjdUTLnjKnKQH6c8tlBSJSbS6giRt
GYIOGIpeVMj8oOTCFmsKL1f+ABg4kI+WM+lZLGlhHTiF2ICF7aIg8bH2DjuFADfqvJJL+qioe2ui
RpcwBLsffho1pG1fJWId7iUhwKP3xAq2c1Ix2nVDpH2c10bXQSooYxLiYKfm8bq+JAByZhvkaJMC
umuAag43bz9hzasjRkSh1sXqTF6B8X44AqdUk21eC989xgtkK/uBHWzm9JK6D5i1SOQfF0LAyt1d
nzEJJr09ANlWyX7tadlvVebgeD16vMOM22idfd5ffllvrw7e5QNBjcDOWXUrc8Zbt7Hr1l0OQoI/
PmWm3SkdBNxIwPf4CmbLOWjaU/VEq1iYdFCJSQfGTCePfol4AIxfZ203iWfLHjXzzKL0GalMTzZM
iKlyJZe0lvQezOX5QxcaXD01sDMOLj38ZvyaN+jHS1uKbHbaTqSohppN0821QZ2HjYEqwmDM16Qt
78atH5P4KGQUNHi19dZ4B8RLnkkyvSCHJX8itJ6D9We0kMAlkce94FTq2zcYLaQ+gorbUikAKbl9
e018mfWjuZ1WZyQSMVxGA25+aHjqH0m/eb/6QV4mbq2srMFz1uJyXvCBXYBrbF3cCXgMtAZXH6Rm
4cLl/ZEbA/p2Y3kZjZtSqnlCJYgLshkJA1Ybopr0wQYMRVhPaEkW2bQXe64a2sJoBzCEwKW67sNR
lTok11AwXRjaar0GFNT7k4R1B6aDni4FRWoeUKJHWcJFIgqISiRCcMCDrYDFDn2FS5Sdw3KV9kDg
1ixYtHtoAhAbfAIEEsFiNU54dFXz7Xfm++kF65pEN4JeLDe+arR41fo78oGQlXNM1+Xuws4mdhux
OQAO4yytXQRZpqpFAg6E5m5qTAuZoMoKgMowBR4yPP21k1yuka+cYYdx5VWilFsk4yP050lQmD4N
2CohbVX0zvWKQGWBh6pZDTuhysOWMgNOPJ70jBjCE1Lnm40OtjSykavOdrMMaSQ5fTa+CQtvOoG8
4VlCURAGFcIW5X0e/fTmgezGtty10agIGUtNGVytpq/dXus6rpBR8ju6lChckLOX87ym7AfdXKh5
yfihOwnp5QVx1hKHQ+1XFMLJyE1rbqS8faXLuspncJSxRSO4W4AORF5d9w3gu10T/KqCoFWslNpC
7pB9r34SJJUolKtZGl6Z7I/xUoq5O22NQT0nsmwPSxqfE0Wgp1oZUA/H5l/3pztN1MQhEn33YBVl
4z9DJUXr58TZNAo5F5k5AKRjMfQ+bDwd4R2dzYzdYMAChCs10SY3Tl+QXp9RkazdREZ4M63NJ5OY
AQH0/WnZHTWu2R+RmBNqJFdt2PlG7WeAs2wHBl15FOGKJQbOl0mPUuz4GOqeyUGOqVHuB1rQkLUS
2mLyJf09itK6fb3YJLY5R3uC/aPvLykw1orvMqE7cfuM/e13t3LCN+NJxL1j+h1lL0lMCwrsOxln
cuSUEFUbnnTMbctnlHfRBslqlvf6/LuAEPdwPhPkIqvGET9zkms/v0/Q9uB+6uX6Uyr2AZRrdtJZ
P0EEXoOJbVzuKCH3f7kdyqHwuVZ80GT6USGcxPqdHbZgLQF+G3G4XGREDPHPajBKxcycVacGrNxK
IirHry9Nrukn5NCajd3QKaMTewVSem/Qv8ZIJ+ytt/uHYthX0QBAP5bRWZ2ncHcJyk34HiYN09To
rccPyxOa7ApbGOOWgamR51NZmvp5dnlHGOUv2PsTWDH4Vdew7YWJoKkn00g76+4uDFdt2YLDnfyD
y3iL/cozq5fArDjGngwQv6FnjwDcrqk3+Gd7+x981vjw0Tgiws4VDgU0aZAR7Ql652P60ZvlLrCV
9k6GWIhOWgaW9j4GW9oeSUiQyyuL6B+4FT7r305bR5Boe6CapkwsDhxCu2INyXcP/Nw2q0Y4UgJE
CwNvToc9HQD2DDqUB6NTdTH4+NHt74++tK0EDOeqK1r5R+RXk/0KhVEGyrr9fsv3NzDqkLDsWyLY
FSgeowevvHPkONbs76MTOVYVz4ZCvCfGzZKGIiqDnlcs/1QO2ISw4u/MzSMTkDEhV2aA6hzlgHwI
v7b7nyEOLJKvI1P6xZtbFEThcZ5K4q6omsviQjScyRk9BqLiTev1OSJPRKzP8ybpyZBwh5Qg8Fz5
nvuNFL+hDac9K7Ys5MVhDVW1pcknL8WX0gUgMEbQAoZlnP0vvl3iPWZokB4StA5E1OzPWP7a7c/l
D860P9GGVVRbEtjT9eXkbiD9vwuX3hNn8CWcu8kzpg8cmel4QfeR0X9ErR+9uQfY8p6Ngo/jFVPR
yH3m1WhLDk97Z2AMFxx/EPHzPc4VA1lgJVYI4RsK1szQ7Pv9aHumXJF5io9KP2rvLFcdpjeviyzJ
9ZAIKBpBRpyYhslkkxSDwiDRu+dNFatSj8lfk9ljEPUusUcDDm3V9WbHtb8FaMUohUItyLE5isuY
kJ2DSSsRoe4RE0TOS2D8jCqT4eDPtFkY+OcVofLbeNAZ/NYhtqd8a5dXOIk49siYDGQ1nEeYY3fB
coLKzQwNiA4NNo5il0DdoiZZXj6rBUdpcO6iLuw1tXSH7SAYFQntDW1lQb9+n00RatVpIz+UxyWu
8ALItndUgK6RTwH1TbwQ8h2uxg8q2kbwOBgle/6sKDNoWqe1kaYhfkycgcJv75wvIPhsJLyj7ZSW
iIwBenyWAHmOCaMEhx1JlCSJDuEsNGPAV+IboWZ0DyaLKiHretBZzc8p37MwNH2Aa3QwyeB3YMOa
c1sLMlYigwCrAFP5iX79bmUDt7Ggswiz1d35M1MSulrC5CQouONDM2pieZOoiZMjdTuPcRvuFxL6
lnULFJTEGnbXsc5ALShae7bOdTvZlorQC+lV0FJXz64kvH5YDG/AdeDdyF5ARyxQYNzRLotHz7fM
FtsRw17q+XM+2VKA5nLd1y8JLjmNpH4xBuVk+hFiHmqoBqbNj+hJrXUR19o51yPKukLha103n4r2
hpF1LBrZYI0KbWQhJdGaihALspg6xWq/NdbL3U/IRZ+bwXMzL3O1SpdEGxNSjaEsJfH77/WAoKD6
xoPQYysyMBT1F/1aCCRfDeFFmb7IL5cIn85NeFc0PAGusb6NBRBFsLqldKyfreSoPKPIYlPJhP9d
le3jKFLEgmCJTtefVXcuUvRbekVO78RyXt99yKBseHfMFU4M/QorqafsviT3+ZR2N20mmiB3j0qQ
FPYlKKxV0UzEDSgDjihx0B6okjlCTEk3HLBuUcYCPJEI/1TVUP4KLTur3f9IFVy3gBzCUkJBk/dg
X4/LQ+nVD3LY+LuNHtnnNIuL9iXnKRSKjzm+t36EpToydWDguFfTFPR5wgupEmGvCrHocn9oi356
kSrNlklODo/VFhyhsy7u5llsJnjEDXDxtlF8U2Z+miKN4vijesQNuBLvCklyhqwzNN/wI/aQvDbR
ilknKV8/Z9ID4gvFpTpYX3xsIllDGktVG8n1owFIH1+2e7Oqc0Y00WVI5nkjAmd+ZdW/GBSiU7aX
gPrOOmxzimOUSlKcfzmyHioKO9CvKlkuxedQ1z7ruzB1kROfqcXHzMWg4OV87VBxx0GslTy4Q1Sa
qLWUDLrvLFskLjy9AKZX4J9EgNgjdttauzxooX8y3tQg6JMWAIVqXRP+o3OnZsv5UYG6o5XmdtvY
BFCbgPe2hQqvnL0Slzki7vgcyMZocSirx8i2CFF17tn3nauQjQT935AvY9HzZGsgkn7OR7kFw/PZ
1kut2O3ommubTXTKBw0b+cjVKGKDk1oYlxYZ28qFVXLKhBo7bE38JLrhEG8eU6V4xQnab239TDNx
Hl93C84Zl5s5Bme4QCDbp/7h5n71wT7Ak3hFAovgC1WkBKOCTwsAHMtV7pjj/Lz32Q9z6ES4t2co
RJIyq/aFC0n5E8BE4rWHulViKMTDk+4xM3VX8ISu1tXZVDUmyN+Eps+r2Bg8Jvoq5BkEAw3UNmuo
6fm16+Xr0AcrrR8XMgJ5Y3YEWwMFfv0qk4jFal2dQCsyttSJsuaXDCKE4nkdeaH7+a/DAbvXFGSo
LcMZEBNwy3KgFJObYrjTS+IfKBY5dZo116emGg4ExLSpB7IYvOgrG+M8tQJICyKus7oNa0vQIjZ5
woDAclhThSeW5bsJIJltcqkioc6pnY4ZmdrvU/mL7A0rHmEsshl8XQu6DKHCrQb2TUvLOe+vB/4z
f/KP5DanEed3EuV6gLu+SzAU2MogmSlC4BZ/aJsgRFVUcxLtjMG2CsSYw0E4eqeLU0ACB8qMyU0V
MmMyYkBTa0bu9zkpYzmVkEPp40iRU6N4Q7UIiA4t+51fMdDiyuJE3NlsIF6tqCR7eWlzBTTFOwbs
r010qpZ95ugZ5h8i9sxtT1ml/lvcjkSCOEiGlteiNKSgzkU09t+qqt+U1VtVMb9256596eEZFk6O
O8aCkIPCw3D7DhN4hpl5qNVuO/h3XzKUjRYD2gMAtcZF+VyhDGYmYr6BjeVx5sUhanK+umCGNJKa
AjGAuty/gcLZW6QFg0jekNEu4DAflcl1k45j2YcEn+BkDhQDCSC6xOnaq659m7CJOwPYXg1hXaqd
FFkEBB4IypYyDFy65lIu6C0iJluB9hNoWOXZOHoHGKszRTxMXSthtzX0cUczphcECHD46TmyF5UF
oqGi2bpGVLPYBirtMabQ5bk2LbKnmegeOrYqjfpjjcmzqeAUs5PN25fWPon6bDoA1Dp+U7LGptP2
exutI3nJcXwhC0qKe6qyX9wLoQAM6+BbGfTAZXUUJZKvPbSidFdJ/PM7UZU052mFNKSAFNcfQzjI
J0LvFiUTnW6GQNm4SftPJ7GKuOA8iFZMLZhgF87v+TduHaBkYRBl0vEwVg+/i1j7UIvdW4b9J1bp
J8MkN7cRma3wWB5GiiF4pARp+IEq0Uz1kqNnmMdXARr8UNScOoQXAqyFIKJq+HUsQnWZhVY0+v3F
hJI6C3DX3BQwlDrDdf8VPNaaARQvg0nmxQ2BfNC4XIA3g+sfFYazB+6RxF5n0qkce1z9e/z7pQom
llMM7zNjWkAP2Neatpb+eyYgfv7z5ZnIQ1VabLp1MyLBI96XVzgoEFZMJly3+bTagEM8ewstpt/j
a+9T8qvtrQLvaJbxA5VnXCszghlhsDBWdVgs0aUxuzIwguyrCr3MfWBSu2XpBKbT+s5+JSCTUfL8
iwZjoajNVCUCL3801b2PA0VpnRqmiuHRDSvMReO1SzjD7nJVEh8mc/HOOPaAZi6bBpCNAsBDyg4B
KyxoyYImNZJggE4lCAOVl4cwC29ws51L9NPkrzNVd63gCjl1ae4ORtUOwxtJ8dzxnL4AiaiLQjcr
h7s20PEHCx7zocT3iyo16pWE2Rak5GIE6ORxkMAObI8HycQpZgzPJQJ1H60S58EVph2lMEhye+5m
uiUqBKfqn8G66oXU/seOS4zwPwFfrn4JoXdckPM4ogwIDJTk56Gg7I7OnaQes3kWMoibDkGdD5iF
04Tx7tZnYXn6Pj+RIpSXVj3V/FgKJvGE53x7wp/6Zrt2bs+4jmCVBNF45nngwZYHyuA7bcXH4HDx
LoCe43KlIT2y06epl99u8jBLIfBc2Nec6Zm4AEkAMQFgLMnVGzIhI9p8kWSBuD4k/VmVrvk+XibF
8pIm2EQutpm2a/qe/yL7F2Hanl1M2OU5W1t+IXbbw5hYylFLQFQCanGsUom9VIUbJTPQNgtr4KVW
/mCZsGwHUVu0tUwb602seNZJA91La2GlC7BEZTz+DDTUCS1UF1a5TbrWh9CkyiqK94f7ZdPO8Ywq
ODpCnkqVeRwBuxxARyuUk4+ZIBj9bHTFDhYSl2g5/gIqDZqdiP0Pxa7iBMhNcjM5y5M30wtFCDkS
nHgfu/t9JoTTkZ/vEOwrzajcrafEUoXIwGFfGGHj2kev0QmnUGtGv+RUdfy9c8vYt+PoD2IbyCzS
+EzviJBAvEBSAEwmksYrC0omQFlocjg9WAEGBp1/ghV5qMMKmNG4wrJIMAIOlif090Ujm90gsTre
kzgJbPlyF9DI2wdLC+02f20aeN7g5zJzxkZnZvS5tmbSPkv/VYwZ1NDr6knNpNSw4IHzT4b3gnHo
o+qkYtQvh1QS1Q7PRjyjiYo/t7NTq6oiW0Wvrxk8/lojqkq27G6y0zdq4hIoXa4cOELiDlj+UpTj
DI5yH4ulDpPs27fKwr1AkYSvKcrB2NDNnJfmy05XfTe07CwkndAVSGA4w5lEL8Eh/uJnWPbksHnW
cvU9hAVe7SVgS4ht5NE0eYfNtPXm56WwKXXqB2ovWV6Ogt2aH2wiHwvMskviYHbJLoQ+4GxXJ+nK
JPzVxVTbp09Idd2JnkFNKkmTMuwDInlQ3SK5wCE5BMSh3omi+NKscjfZmOj6e8SEP1OsmDit3p9n
MuKuVCSr6CMY6GhWjWWJHdp9VfsGSe5UEhMgkypZf0rPe5nKfOOeoErcEUGt8XAtaCy5JwtPYv08
AIWlubQtq7/uXxYlC/wPgFlaxTHYRkT2BrMYbj3Q8FLmhylfhweFU8I+ppNUj1gjc1gc1iK7TSup
3e+mDz6NEmucOEYy1ZW6XUgDmPmUEDqAlx2RkOrYcxWKfIjZVO92imSXtxexkTDi4hjkR5EqHS/u
T20/ZtDSqoccYRNP57JQXpD0oO90z+B6uVpMq9rJW+7HIp2nuRv5iAMMzda1Tv2gGAJtXRfW0Pw2
49PdFMXxKoHUjakGgng5gHCGq9Na9+gF7xiORGYDicGntDes9ea0XONURHoEhfbft+cBsFpoJ835
oH2BvU/jHsyOo71vVMjSWB/SK1tEwyjD4KDpvcmGjT6j1KI7wM3IWlxpuglOFbxop/q2PJ6hscY6
hL+yZou8ygEktJBHmehYrGccmFQy00Ze1imon3PyEWufDw77mKw+8QOZljvo3ZinKpRUhSDEcsu3
RVbiD8YZS84QwzS76zEx8PxUiK7plAwAyjnLErqYymw39OtNP9AhjMfdH54NZC+z9u6AQnrtCl0X
3IgHxVFgJbyJHJymJ28c0WnCLBl7P9tWlE5LmEAD/x11+8jAa4I16YEUsoTnYOrDfhtITQYMNRDt
OKhKBUVIkh5+UtGs6BiFbekakwz+WmepTkvQ/5haOn9YFK+wZS4aQiNKAEzu786PzZeKlEZw/nvH
l4kowYT5uCUJIlQUv0gvEnKIJjZSjBFxkw5FtA4rMFH8ry2PjHhKwQZ+v6QFBXN3JAVhJnC/V1fZ
oktpvD3r1R+8wYwQKi06YjmDyCOarPxmTWcMP6jpFK1aeg2qBuGVDq0m2i7SM26lCqz+KNFiiwMa
cEYBJ8Nlk/xTlM+Wcd9WLD/x3BIhtZeRM7aNq3SYQHicCexzWX3pq5lfL8ZfFWKrBOd61I29N6hu
hFanJ1Q7EkaPY2ltmzADP+KDAsxBQKWs+aHm1KG7rlTzRPPyyWV352l93DcxUH2g0TqXcYw+zB7o
+V0tCTCsvN/lGtIfkELcnlwsXtInLOIhexwbL+CQuudupTLJdv829KEmG2DSPiUfmklji2mova3z
WLHXsBaK5PZsSlKUJrkNL/gSE6YYnJQjnTfatWdX4xa8J7gim6iRJXwyViLVIMNphuKrCE37KNzh
Ymvu5eGPQ7qjJ8msPjRmvz6XP0diJ/gdMdLYuc2oMUYMjNYYA/3/QJVILEQzPuk7HaKJWBG/MCEc
2G2NOhdxMxi/HQ+W+uEmdQz1ZhNOx/EbXkctzBVPD/pQiUnNCxQ2rBa4pfO8Mo8nHVPDt+ZozIu9
sdAHAlrPQ/4PXgpedS0tz7m92+QoeSo6PtTHQa4CTh0B9b1vtPofO45pE9dkzOlnHcO6w4lZSBBN
1ZujDGaMnphtzUjUOMzfVRd63LahqTj6NrlsBWwELgDuXObE5+yXTqnTe1S1yhTUKSgsMWMo2vrc
KGu2Na69fGUXHpJ3EA5yFPjWBEwJbkogCsS/X73RKwIcYzx8nkanp7WEHVV1KD81XLnSDX5VpOE2
aggMk9EAhD4Dz4bhvV5wgbPSH+ksoIjfvY0PuTXPXaCl3PngDm+/E+/x6OwPy9yWE3gnpxOk2mtU
vCnnv6fCnLFqCJeEYP3HTVT/aUKMhWlknH1sm7WCF+Z/rNgH/ZVulriEQVpDFBwti2+Ps5TYsIoC
8a4k0+fP/3lBxn6PIyqIk8FxoL4DFdEAAVJmLZvViRtqC7bj2nYi9d7eNaYqFy40KJqeFOcl2Un9
FsPyUVHVFfHBt8Y+rZD1coiZ1MV0z8T/4eaaWGPYtE1nu+iMSSjZJtgfVJkqNyzo/Fhk2/aFTrED
+TM9DV3De4tFoW+Aa4TwAp0XnhSiEXs3lZr0NdIO7CzFWxR9AFQS6w/r3iF4XCTLTSia3l+S+Fcx
F/NHkylp9RgCc0Zp4HGTdH5GlifI3iTETNpPP9Jk/yd8QRcwRJfUx/VymFuqWala6N61A6TNfKk1
kPqs/pmb5TciQLr7lA9qoycxCmRlSGs7XYBLxI+no2e8lMfhPSOjFPYKu1Ho9QBVMDJua4Us1SMe
dLDcJJwyA1JQjCtXnCr+GpCCB8f/isqUTG8xHGtI3cUvA0Fu4GvPyEsRTCR4rLkBE0KirJLi4bhr
wyEQAVDZZecg6OKUEEc7vzJPfQiktkatUCG2xwoZ13iZZ2R3U775gYhhYYMBW8dgeCZrAHUIBiq4
b2pK+SSv9+CnJMNbp/d3ZtJ2/mo7ntK+NhjtJA+pGAwiRc4DKyH2H7vLAu3kuyPUcSMoIxmDxKhK
l/4jYKYEUkkyd2Ivt/Iccl7wg/myCoDzd1NDN79DMQ3Bf7qjbX0UnZlWmhx6lElDrVVZa5yUaSfu
rSHeflPbGehcNcQEmbVu/o+v07+iUX4I5rJwU1WqU8E4/M4v2RmIXBg5MZNp4qLw/OHdFmfHoOlS
XXZULxQxS45k7UO1m4drTDExMRYnpCgLgrjr/Q5tM4VdnAQQCU365IMWoBb97qAidisLdKADEIMa
p7r1dKp/VQNG6j8rwTpMd/zFJ90HSZSynrlyeTF8sIYJyOvTajaZvflbLAxgFgFODvfdN1oC2pM7
JaLBbHynkXcfA+r8WOjmeLSI7W/iNvsFVsasoXCv+hVuDTaalq2tHUIatCau11F4dw1E6k/BIFr6
tlge5LTff3bQWYxk7Q0AVO4a+rkS4NBpBb0HLNYhIx5JYrNRvIJpwN2EB+K+08WxeihJhPnB4E/o
eQdwgJ4qNm8mjMMzs4zGU+OX8dC6zjsOVAolALKNwlD8erv91SoveqVtU48v/cTwO00vB2j0HM6K
ndbgdacP7biaXE6Ng0F22vW0BHQY5HHaGZCGx8zTz1rEYyVav4XRWdyS+17sS8pEW3K2wIxq4oZF
xq5nI4dJBGus/5O3AiQ/yLE3aiSY2fGdo0p+NvlxKfo7zWsDM+xK1gJqp3kE9Ucax86fvvSMDjVA
72OZhI5PDox8kbQ0PMpEhUWm630t6bIsGDU9zDKFGs1d4RhFVtSDbZM9NIGex4HLYaXNQEbKArN7
vt5lg0gAbtZb4Agbuqxeyf1bC6uYpKnqCe5s0YVIqCS+wU+gz6Xn0uktIorfCRCyLTeV+OgM2DqS
rJZv0A+bey9+jWEQuLH1rioHY8/lUsnrCaGRZIYivCAIfdKRz3llGAIcBfAZn6uNniQPNkyA2dU7
f8ZjtJMXyHV+9iKkaWWyOkiQ61ZuNd5mxou1nUtuqHQ9aJwavviF/wB1hSiLUX/USeziHMM3dN8h
GgF6lSb4tZWVTmwAxiX5lS8uTQ59KNbhbh76xmTy6dzaEcl0jFYXyNBCBc2cOoNEkAp7PI88HGIc
Sb6L8GtreJ2NAHm1twLt1JFQzPz+J1DUQs5QvIl3NgHYin1hUAOVVlvkztq0O29Saf6uUPUnkqFK
RgguOSfEdIruFAek8xXUMXGifTtEAXmYabRtjUnKxFaySs68rWkatAaAOwR+EKNgA65p+s0vyPPJ
+DweoToe9xke1UxqjBv8waenIr7HsLB7TeWEGdYoPBzcasJfalHDG5f3ASfjXIjLIscxbXpyxNAY
N2ZjXPAKAZrLofQDNzfWqQvGr8QyWJSf5o5C/QvP6g7ocwpf6P4gubLPR6rLEE/1ZLIlNwufnVyx
hDYI/xMsaEIbNPhqDtxsZ45jwonRFv8NA1GTVEQyX4U8aobwPfLrW+XnqjMtRFnTtYIJogqESO60
pmntN77cTjUZlgIMS2GFk04jOC+32uMA4Cy3CVZnGQAcaSnvezRMjUGxN2pXnq+NG5h4DXsDFV3M
tSdwn+hMKxjvZ/RcwsopSnXtpWpb547G/T3HmK3CAvpvpMg7ia8DCnUMiQH9RInoMTFmunEJS25m
Zh2iMZ84peLmNAEMT0Ck2OFiylhmI8KF1I1gjrXsJVNS6AH+XLSWGmdWUnBinCzpGuWjkkz3oh0z
DP6eQGA9MoO5CUEykFv8b6V+V8arm0pOqP3CzbETFPTX8/8h716rQvdv0esTeVLhh7YfkNe+JRBj
/nZ/zElKeJOWqzPIGeVbuzW0v1TEMlyidH8xC+kIhvAckG3fs+7tRXNAv2k4+PwYdEQLdOcowJdn
oYVN+6avjJ9jEegxwVA29bB+shhdpQ2+PybpQfDblOr7Tf0qyox2c9nU3DrglhnJv9P7agBHWm4L
NtsFUGn+x3T/CQShaA2m2QRI1ZK1oc+1H/7HMfn02vsQczJlE0iq5Lq+UBe/aZXKQQi4Jdah1CAh
qXvTmxhk0t+vqrlqD4H90RRH1TjfMVUCqp0dJPP96nUV/tJPcPuVcynGlFTNIFZXRO6BwqFEnqco
2W4maFdjKtttEqcVTBtKumJS5Xx6iCIKKexbiBEjehKz+yTUE7swFB8VS6LEEGfdlqJOkC0bPsLZ
7ejhp1tS9siV2kRrXjvWjqZojg2Fs975YbPatitGET2SO4bdOKOJGDn80twHF1afMhCYfWjVKfM2
lOON3Ed7+2QCPU7L1S3/H/ksy3+wF+qCzLrv8xWhL6c9S0/jQ8xg92kdjOA9dWT1FqJ+s2gqhVCz
GSZ37RdIF7F/dF27oTkaI2xgjw40wbJqWXbdJFxvymjqvDL/+WC5M0Brtk6A1IhczRVCykFB/TDx
NmOt1MYWkWGh7Zk6g6ZFhvSGDOi44C+KZi29nNFSIPsjArDKOhbwFaEiQCGVhobbHg7i/rLMIKG8
gwrjL2PqaVdqY0JMmfi6DjIne/9rCuNq56ujpjXb1odb1yECutKSQ7xn2HjZ1kP+CGznS1OVz+eX
gAyxAaFYHaJsVRo7zZ10gWXqX3I07WJ83dTA0/c6ka2Zhq18c6SqR5fTo1NJ8gkhkSRXaMVwq3Am
HAqUe3bNpycoBHsW2jH0/eAfy82b9Bnl9hTpH62fa+kmYNS73wHnn83hXIxOz2IET7pHUjwX6rYu
Rcdyb+3y71XTACIJLVKXc6ft1dgf/qLKEqaz4p5dGX2KNn8hk6qWpgi1xz5Ki4twBkO1tMqj0MEU
aY85+lqRpPlPSf2r3XShP2uFixsCz+/vRevptWSubetcUbU84aRCnGFI38PdMkbigCwgSzixRRpp
tbgU+0Vu28D3PxUWoYRtNRMPCTSfWjlriTD4h4WBktY+NV7Sdw+8FiUYGnZkANZmiPZyfm1/7eZe
RQZ2XVxK2T1mlp0F5MyRAXZ0R8RZBywf3HwCCKszdAH+3+G/AdCzwjuT0Ad1GGEUfvtko9vrkHoZ
MbrP4JUF0xPMHV62kWyRfn5DFMFMYdYgV6qOyCEjPxvVo0sXVpmWC03lfZl6Y8u76Vtxd3wvdDUz
UCvAFqIHajqqy4nkuIqq9rIM0I4bu02P7NpQy8B+5NbZU2d9r/MoWgmJWmUGV8RkRtesuLyJmer2
xzhnuotjjmvNwUcXVWM0Ma5Rg5o+1vKqPysmuhmHE7y9MUFRvjtDz9bflxOFBeFbL4CVtZT+0+7X
RTAcGPs7dEuHbXTRTEMKzPLeW1mk2ZklE4yB+Q9ccdKWYRAGvWigoAkirXBTTB+7W1x3mmBNlsuq
clq2hVhvWVcgaYErtX7Qr4IJ8rPZgaMf+qZVEYd4IcUZ0BMMZgWAHEkxV5fAEnEoANUj/nOBDKaJ
0cgBUUBIRyTOnGJs9MBKyoMc25uLdNvHNg6zTWyygThmM19jsrO0jXKAKC98tPHDom4SfzQls77n
hPfcHuSqxbux7vWZ8gjsVc1uomb9/f97WBPYZY+JpWW9OuitPCh6ZVeqmNOTtqAQZCfVQihFB2x3
CGRUIP179torRUp+R5s3b1yKZjyKzayyOmTYi4+lEU0iyCsuYXVoFseFV1x+1P5HtBvinyHouL2P
3wl0+v0xQG04JtKCtdJ42SivzRgHTff5muqq1Oz6639uB6UF6dAYWKCGytGJ39Gg+6IgxbzPShJU
h6s2+5bEoT8SpRYseP7yGQafUG/wjdAvBjdOCTBz0hb3JYh2Oizl56DiPWnCHoDm3Z9b/mEaM1YZ
k52wwgUYvWpzdgyolioB1HeydpvMMwFxBj0cV4y+c6jB38IroXUy1r5JjZKNMkjzJ1rXaoBFViG4
THNx9Dyv+LR7O89t7y0CzVjjMMrFiPNOBqQPWcvVg4KWlzySM3FVnRtctQAfdvDkRZpejIEJ9QiO
o2pXb75w9L0tBssp+D2Vjo11yoFjDezW3pZ6X9FIfUa1iMfqXzKIohZaEzo0AswZXqGx9MRp1h2Y
scb0K0ko1szHpKSMVWbFADdj8RTP5I2AZZn96mNforI4URxoRQX9AS1F5bgtJImwXGEzyCFMbHJP
gGa86tA1ClqTr/KzPvirSs7PIYAlB0BfTl5mwVFT0kwH12SvKmuyzVpm9iBpX5UKcAtkLqo9SlxZ
giiIfrDCFmK2Q/yUYzr3ek61bWWmO8KyXX4Oj0oTRbDBttcQQAvzSbVQMYxs45/09aLfWfW7DKIz
RGGbCBwMUTgwXLXhRNHmZAfL6cqZDoTWH4lAYKmzcxrPBLmymhEzys54Heb4avqOOWdOVFBFadHk
8E6NhVV74jwfeNzOaL7yHMTpGtpOaOBeSAebZLlOsSQDfb1g0Mk5cWlYuJUMX4fYwpPNErQh6xD/
z1pw5wJ3A+F6Sih229ZcKVBeI5aoG8IpNRKC7onlaQ/mLy01B/TyEfz5C2ZiCzBZ0oN6E9Vk3wK8
iaTjeYe7oJ/pqNNMen9YLlV5neXUDQMd7eDplyvDyaem45GU5M7fmblf5CHR0G8QBCxrQf0eMPZB
ssxUjmgfHfcFjBGgzgyVuNacDr7rs0+fzsqe+7Z58ftGKC7DMmBtcFvI7ZU7j/RYANsg8smxwvgC
TDARNJvn1KD7f6nGdOaKOSwsW5+fhqewBbaSYDobazhdZpqvvsiquZQM4VRKQwxmhKAxnnH3iLe8
WfE7ctMWzC2DMFRmHwdmUoKSX2tJnG0BJqfHGafaOwUc7z5EHG/WNfTmQ2Wie3rHIXM7TQPFMKEi
JdJFxessrrR9R0+rpcYVohSv/0XacmeGUp9Rw8ZjmYwWyn6Q4u90BALirNiegrwj28kw9NLSzY1X
6YKCXz6UXH9UISjj6vE6wAeFpyieu/rbbOTL7Azqu3cLIVNrczzwmcySWVrxpVaJzlZrymdvA9LF
PJsq5U+9Riyiy4HSc20ssaZGO3Iyl0/n8yWM25InMM5dzPK3z3guHYp+g2dyNMSa3hnfABPBgCnb
EWBoUmjUq59IjhWQ7iHlr80CAXSCxHTvrNPkwXPAl381SKZPI2Qs69q+DkLEGZSD0tDbmsbYHdbw
8W5qqraBkylDHo3Dawcz+e2V5X9RTb7cEiQ7xK+GzaV4Nhp1BScUbx+vEGZAytakM42tqK90UyL1
fvYKeSZw39UgI+KWsMpBR4wkZBUsKfYeZlqLC43SruSkOyOTad98J310V6cmn5RCMdO4+HT8f1ZG
8nQzsGFriQe7oZ0r9nBUXfaBSu59uG+CdY8F8mPfsRKqTgwFQvkpVZWQggFxi1EZMRtinDz1i2oB
8atMMrdlaCWe4subRAkENR9+8kZuCbm0C9dipwfpQxjoGSJmTcPNqBC0+fEwvyuSWtdX0EMH2/X6
Y36lsrke3BUJBum0SIwqa2yr2uvjYj5B7iMZQoYBTkTNGUbFNhwE2yupH54FmDWT3mwxsKiapoaJ
0Q1vpQb5MvjrzbV1frFHft5E5V92Cw1sZQTLNAdyL+rR6ApL87pxm91IVG1RvXavE+oPiWi3li1p
w5vKnEKYE9TI4Ug7xLGYc/ca84sjudQozjcSXH7FPVB+xQ6VIP6Eb6wNXS7QLDOlhLnj9iAwVpXP
0k17xxWyAddOmEUo3f8j+pYSpn9eJ4aZtFfZS+S94RAgRixPkgiu2nCRNVKlKkxX/SqtnimnhO3e
HVtKHmrHSI+vuSJPZOQzAbhJT+DQT+qDo9N71SPq0T9pKGTKFa/Shq4n8aW7Yk4yjGb2UMx2UjZx
efCYo7wFwXnPnDqnseb8SnkufI6G/C88fYz/nMalMwlzZFLUvp/usGTlwuLWY6Jq8puRTo6Z47w2
UnBpXSmksiFWSytZYTuM7KcaOwrMIFhNEt4w6I8vNyL+byEFTsexR17PJx+quH9RF0nSaH27Q5bE
VIdgNajc/0sFQUoU8fUX+8eoWx0nhVkSv2EenPueS8x1fslxUDmajmsb/69TP02VHRRtoo7VbXFv
JkhpcrvhaYg+G2dpKz0wZhdpVrSeo48Tblde2JAY/6ATgBN+yWiXxfjvMxGV6WkycF3CjaVcNeHM
cAoh0TAkC1fx40g0jDpS/Z8u2BZbrtPramrx7SFMtIMzkcvw1O8VR+ahoVep8DBA7/RouRlqx9VB
59xj2p0c48rVDm1GMsHwZWlXk75USt6NX6Bx7ipImzPeT1bwL5cHy3lIFiIOP9Hr/7/I3oWXCusO
OmBoFNv5qPk7jrLmgkvU86NNfJfafpLIv6+Ah7/C72gRguQ4faG5YQG05UOvfqk8Lg6xU8ndd/lM
rc77CXN32mwSzBgwMwGRfzoohEJJqnDCWaFFmt96hGOC4FSzaB5DSm+xePp4Rv472pWcnCMUoRln
qf+FHdKmgLDTNxV6+clos3tUwpeTJByxjVF5sALcnTyoyJz1DzB8n1RmdGGbM9QibRI48SFAmYic
PnFTqJzyLPRf7rvBhnpIHldryjO6jhUj9jYYWEsywkxfDhopNq+N4L+tTLPg0N2B3yOaMR0qToQH
9Xi6VXSSsvmBxEiQyLNLqf+EQdwRo66AmH+WLYSF1UjW17ZyUOvCRWB5zTAwu10soo1A1Xyn7h43
WrZyUMiAbiGfqdqOpMH7U7G/KfLC85PUGokMk9ojN0cYExxoE70rPKYOlAU8kYR5bMsRZvrIeSNR
/wi7dkCjtnkYJxDEAReOZ8BiyVdTFn0Ve58wM4bdpHgjAWRbOe/+LvfCwKJuirVNebmYn7G1UaEh
ZB1UNFBljXciHEZh+uhp2f9TBr2pKUjAl/ycbfELl3Oayo6sAO+GIuKnwWntEBBVudMX5FrIrLLZ
YS+gznFV/vURmXAw+XDPdZ6s2c8yaS6ZJ5uLcs9Q6HWZq88YqCMSzUeCOfpLx6IXW9Zh2oIYTrox
kT7oljvggmjOaKHptTPbOmPBk4qO5xR17FAgwyRPSiNVmiwFofk6OnMpQZoUxWVmiEcvJIRQYb39
SClpOg5HdCwJBioIid/4GKb592cMkTcLaG9QAvKJRBqhGUpW7oCdRjJ+5/s62pTGBGnW+LSAJJzI
p8751VLVfBCAL7X0heAzu9UTzHNAi0dTout1qOLOmuYomFoLbnSwQo+vOYp0EvoGAxJR4ALMYm5B
k1S3OwlcBL+jPPQJpwUqNWeGXAUYO1pfPvmdSawKGVfCsOJg5rWJvYdt8am2S/a0eNktrVX7K56Y
pD5wkicYCC+ST/U+yH9/cve7IaEWaVZEt95uKWwrEsykVP3FSSZ3sS1rJg5DP44NRK6TtqhT7IKL
A24yqNmsMfEFc6b6Sl9r+ehu87loYpNpFcr8YGAQR5T88ySce1KXRUMjrCUkgigbh6GlXmEy30n9
dQFSuHh69V3DHdX+Es8QwF+Iy1665dzWbTaKIEhHFad5YBaLwoGni88OYuH2OGkMTEDPzeN0vhHT
h11LKFZxHd7duKvT8mSljeGh9q0lo3IciWeQLbqdZXAHDyjG+Kmibo3oKa9rWqsRQeyZCKWC8fh0
xBBDJgZ+AeJTydHX2F6QZjaPa5Pdgvglyt15I6U13XMhAuPjp118RQlVYbUER0p8zNSCZoKe4kVW
e13yDY2ZUD/Ju3oF+My53Kjy/Pf5B/zkIv+zwRWDR0/g72W83WaMsVwSNQ1Z05PvzWsxC+xViNIF
4WvpMON2gq/ns7TkxHXHKvdSIYs9dYtaSA9gucwIpBWwgSQZe1BwQuUbLRxIVfKeHR1mg9WScYGH
/50RYiOSvE3x14pdTmqIVRaiMQjFhWhf4w+uO0OUbwOY61ULkWMdotjluCjEd3RFArtVk3oYHEuN
K9ZR5aLG/75eYoCZNYMuUXICAF9PqSSmT8NBrBVuL2CPJnHzOApTriJqEji57EzgtxoFqmFmD8xn
rpkxnAmw6e/H4dnlIv+NWvSHCOywP+/A9nJtZEdVt8r8lo/70jwx9q7Nj4NLbMQzvUAElatyaFKl
dQqCi7hitfn5tFwiILjGcHAHNWQCdHEv0erBZc6UxumQwF/WUD4OWJQCw2l8L2o7t477IpCVHwyc
STNcKJGsKvL9flycSUrtEr/hUGwLQeZhIpdTYznMAFn4+MZ7q8sDjw4NWpVcAvcZYmybLucrP8Zc
MBT+/sqQlJ/4RaEo2vuUc+Q1J01dJ3FfRignU+m2aLTkE8Rul6dqtCKgce96gJlN5tVqrkc7jIlA
Cs276amW3bwWpd26fxSHiD4PSUbgPljeKXHvahPXSkG4jb9Z6jNvDz5u+RgP1nDwJM/UhOjFyhr/
b7/I6y/Ydu1+B7GpSD2th22BFSjV/mvNNzjhY0jCX8J329f0BD5bZgm2oy7kh4p28kmdMxcHkfYM
L2VPc+2ENUfNerBNVvfQla5YbMQI29/xlHXol3eTOMg+EbQ1UTqFmvZCR0Vp9fyQZrH9CV9k0itS
lhEZ7+MMkx5KafhrJ3jZDbS2zJivnZBODfyBaB6GkpuklNgF8uouD8GnG6CYQ7b332x2JsGWDHxn
T5+vneRa/BJ91grsBaRkjbCS7nrTBrvgqMkTAPvTq4+YKGsviJk4uWOF4lx9Q6kiKmXQmS9tZBFP
0JAeCAwGHZtbPp8fHI9SptsX8DHhykyRaDtFpyN4kr5urY/7nEoaxD72p8S6Hdc4HZM00DOwdYmX
QqFEBofxi0+k0eurmZM2wMU276l2jIRsRyI6fnhDdtfHKWubM8jh2GPIHNd6zxOEMbNs2VHe+YsN
ZwodNtadlAmQkov73VdwUnc2jkwhG8dDwVkn/SH6fgmj9kv06b1KJbOMSAyDEIgZQrbwATKS9NxE
/oDfw6Ev2kWug5eVdmpIpwusMDw/FbdnRG28E2UcyR6IIztDv9Z+5AJlERcd2tO7te4JXieewF8A
qTtuFawT2PNExDMDL206Q5rng1IM5HG0kbYZk0OxQBhZrNWvyR64IMNcrhqAQH64uBiS8qMF/1/5
mCKxPIGhqS0gOJCTCjqvwqWYdgol0QLYG3T1SHFT0tgnfA1oKboOhpH+IGxGnB5A5xehDwE/cqc5
VPpmrPFfr33yyP/7vx9BZwYyeaOY3ADvNtn/PlUJWoh5GDy+K5tvWgRiCdTHu0tmtR2s4tMReb0J
hKedO3ixYk9ExTCsCUVncwJj5BLXFxx1Vz8mk6S6uQlhHxlKGhzHOGRHZfeuEJlBV643C4NkxfB9
8h/fyeihktdXY0ZiszbWIvSc4Jsp8QH3H+SLJS7n4pa5pStLWxLZwifXiqOmyyu9E/SIagiV5dWw
hoo7rvqVsYzm/FgkstXHaB5hlUY+9eavMeG17ZwdgA17bEhanUgGziXX6Wslh1GCxEB7c0nlIV85
ueqkD21vqLQHa+VvDm2vXv93Vo2qOwY4MDQBJruuiq7yIAUNM2K9HEzWqDonDyLdIM5pa3RDh55Q
HTFuzDP66oZVWRxw1TJTTbcPM5AvIyhwfbnP979Wi5WgDalStHSGnpo1cRekO7+Rt72/o3I1L0B7
9F+gtgI7kcXYdZwVJpncVs81ykEYyT4mzH5Tw61HfLQi+xE7S10yS7zLwMdmO3jttdnfepoqh0vN
29Csd60/mecB64D/1IG0T30q/Ot2woIdLEHln14GF8Eq1XKLEthPOw/LCsn4NFCb/zZF3e84Yke6
d1iFODJDvD9Zp9d2NUWGDnVLMgDlNXmfmqGfMPpdAT/ehubdvV5L46nSSBdgy2/AKcqDnpgB9OxV
YmCJo0gXrCwyvZI3IqSrU4vT7935aGNLW9gbEl/rn0/71rf8OPPip84RITszlljp7WB/fVW+bzor
VJAI8mlxh784yXY314tv5Vsi/u5DI0c5XdGewQiQC2w52+eYbMenYmNUshoKeNX3Bz0lCwst35uG
pMzDxO/HpcqosdaSPuxZUTx0P63wgotMKnBwD9zH9nYG834br6N+Ui/vUq+2RMJ2ZB/MVzu11i7R
es8cX99jm1d+c4SvFi45mnvNNG5WrrbiUS8eJkneKiFEZNpXaUqMYr36EnUCaEzxhkwmFtq8HwQv
TinLv1efUAx7q1OrogrV0lq7jtSkwLSnr++h/V/iLdXTM/qCXKoT3+LC2+pN6OzHFlqoP4unQY5Y
bPyZNgpb79ilc7e1u+E6JTqjFlP94VU7TSPYWUeKNc+6+02gCqr4w3bx8ButGBgeb+6rhitt3tmO
9ycWT/rmpwnDU0WwWtphVczqs1EYdUQPWL90zyOsRZEWnZ98GCcE45XB7wMzqeBCHlosp4MhK2P4
xJXvZoJ0Ujfrcf1+UPh4CX88L8cqVEhYMJDf5c+V/mpmbeVnqxSHwByvh57uJpxkeB87225u3/l+
lV9hTJEEVEv75+8yguHyijrB5fekT13AHDAueLQe2sfG5I19xkxC54wWg4oUImIp78CE4MDa4D7e
we6BxpXwpqpW4eimjq2zEZa3bsGHLpbI6ZPBqRm9cJyL/apM/6G8VEoEG3bwDY+eLTcRFNSnBBYu
iV9eu5AQcu2uJ82uMb8u3Ig0NsS/I00MUWXefkDeww05+QyoqaYdhn7xAuLUgRWXLkQDoIEsqSpn
9L/YOXJv5H2ZOEp6xB1kcFfpL0c7qkSmwu9SixILZIuzY5S+hEY3fbJGMZ1Y9nq+6vScV4zYI3QT
5aUGPwYtKog9kUUTFHZADhoYUzUFxEiZKhOOWCafi9pVHXGPIFmlt60WCb+rbHXUc+D3pTmisdud
Mkh0h4HkF56SAhSYLa6cXdQPhVEXqyO3tGZvPSfuaa1pCOIelnWsxu6CIRxC9IGnUE+/l25O+UPS
y1oTK9XlVDCmbzArNacDj6f9qcICIuIrYEV6zq/AoZRdfXugO2MseXWJGBTCP/R+LLndxGn4IHcY
Q0ueAvOAlknKlMZFtbiAFcfPcl7bx5WLzA7gqnVegEVbGzVFxOQZop+13Y7+nGNEnnSpJUmss4xR
e0NZ2HwB215kIygCu6YxCt00gTHAMZ1/BmajuZKU/aSC2Xg+OSv8mgFfyT6pPp2wEC9lta7gYvIl
BmQza/Z57nHsj8VvC5nCY4iI3qUpTaJVvSxwgSsiA59IodX1Bgxz86F7boOKFYgHxSLCLUqi2B1e
WU3VqO7uWPAFwKgpAOv8Yqk0XJnafilmT4juSLn/31Uf5zV/6BT5a4qfj3w/X8bJe7XQt/nwhdEN
zCyEOWqGBV9hI3IUWSz/RIc1hqCjQH08E3Sn4kh2lpd6OteEuzZXRA6uFsi9V72wa8NSm8Nc0Rak
YBpYsIWW8AjR+jbrEZ5T19tN//vIwt+A6Bj5bvRqk6SZLWiioj4wg3QL//2Yi2cRnSiyMvaDYv/3
NoBR2G46t6LurCKSfV9xGQXCpJ4x/USRMdLBO+pU5tr+5fkNN089IOy1GW1KATGOmcXT4cqDvg3g
GMcfUpRzkWa5hYRIf3ZnUlzVWbvdC6NU2Nbp1u9I9stpu8aeRTLNlYHLiehKrauCW6Ses8bZZiYK
u45BIwym0I5PDgukmXsy8NQUM7DvZdHBjOjTaBsps214j/9zfxVt0QoIoe02bB7emB+G3QpTjqRs
myDznoEeA/wykAHH2qcZCK2Xh72/d0gCsyywdGdT6lznARNOz6ECrNUPuByA4kqtwjPtX7sBGzO9
ZtJ0vNd2t47cIFdFfpen1fCJRiyxHmsFOIR+YLZMEgcbqL+KFbqdV5gjdXNa2nus7HEyYc+5aRMw
SzgI1v5fAt5b24XOJs88nOVxI2J8bTzb7TT4W5PrAJEh1Blln1Olxm+Mw2upNvDPriC5FmERET77
lAhTjUnKmVaooBAJ/axwNPKKnnfnMS5JkaYWshc+9nGtL/AAvRXPP9DoyMz+v5kycfsJoZaAqf4Q
XKER0aheVjjE9WzumBf7V33Q7J9NdceQ8QWN2XlxPrNXfv5P+Ma/yENSXfCE2oqPgEgJh55msMW+
Vq2VmPhG9wbCa8jQvCCRp8CjJ+xlhUAJ4UQxidXS3mnT2N8T+k7p63fXctOWN5BC8pV/mA4EWcZ9
l+Mkztee14TdpEtrouMXHIitxCVQRz31dlTm1vXfUJhUrNghiXG1bBPdpPvpltdBgSrq/97cZ4xN
WRLldxJ9/O3IQPBxOdqQ1wzhhVhzYuiteGqcndJiZDbuckcjsK/fMZ0iWjdt+q1JCeaFAZzAwdWb
zfyNn2cGLLW7UFV4zJpM5p8LyrSGwxDBKRymEVKceBTK3hmVHn0RWlQrMkgjATPh178QTcyPXF8X
l23eGU+iIEgxF9716O9k09zx+E0OIViWbhU4zzjkQCb3/XHXY364C2jIPoOup6GOS0hEU6vzQLKp
RM4fKKELuEh1s0MZyvgCWWM+RZmCYgJYW0RKX4corvFgPQKcLrp4ySpEmeL9Nz+O8NT+MA1XhNno
SjvAIIxsdVZfhf4i6d+edisoRumBq2nIo00uPQ/UbNBm7L969bWvG0IHVoohUPQxJiymzzIwijNE
FhDu4XmBk3cO91i5XK4DVXCTclNFXRPkLJSZUlLkWM+L7+wu/rT+eFqJvUV/maOIM89KYB7EPBHb
7zjV6op46pBk3IMIyKJTDeX5CrCGWqJRVTOkAtBNLcusUT8G944KvndJYLt4OCgAccMvkDlZzqXA
xRpuBfvz5XbgXHAtdNatkE3kuEO23dL4cIAkLA+9RJ3nZ3r9rgwC9asTbCUnow/t5NPifeGelfAs
49V52lJikGkH1wEijs+oV/amMCWhlTW2quoOukrUasYrEVUlK1nJadjNFpfcLHTjiEdCnvx161zv
oDdoONOOLu14GEeNN6O6bW792lIkRYHSeghDi7vuvGhuBZlenNx+9KbdqH3yJ0hX+RtMyb2L6G/j
IMpEwKkUM6gWxpnFFDeNRLxsTU3dhrdYM2/5Pi2BILmJ8O2KEXe78Lvak7spIMtACkaE8R7bQ/C8
KLQjw05q2n8/VUjz/+PY7FmulHh5pyA8PTEbiqFocsI8KJRx6ZSKgMQOme0ZxkLa6SnSgXLjbHEB
hMB5sbxDHh5RYj1tyma6Gjsc0VkwJJnvi3v1hCAsaEmEaDHIPYR5ZV7DajKewjbZk0orRc2jEk8T
y//GrwX8VFtypGi3ii2bz6m198mJNJoEWS0yIo+y7KshWRhnacU1dktB5nn+Kykrh0rUM+SNUuOj
u5OCb8RdcaSWhjsxz3ccThUWMb9X9BaCSVuuH9UaEutu1fFwjCSfxsQ5YTL36ANYnX86cK5KBN1p
SBVieo+TxyLfpkreziKzfTEnr1oRANIDQeoo2G7DrK7fkLsbsUCO7oXYRD3FlHmcj/FU6lEIVifs
K+60U/Rzf4rwHJz0gQIdDocygLw/RFPHhChFn9MxawKoj9XtgEF6ucUmuRoG/Nme0JrvNe6iJIxq
noYAgoVnOKr00nKCAhiLxm9SPt2L4U0pa/whI/RhSSQ3pYChsm5BB8a10ZSmzUeatiP7aweCzhI7
N2yhl5lRy3gL4jrSTylwFrp9LCkehLxPl2uqP+bcU9qAPOz2QQUyOgJVgzTJHlbuiAnJ+0frp+6P
FkaAsM4Wg7SXztyM56CSRu4EPtP9BMREHA6gQg/6WW6kP8mMJGLttcaqqXGX1/N8/jFs03lKWtha
Gf1j0+eqJ5r/LES4OspT107aXkzkKVJisPLcQC1EHqSDGiEu6iN2l5nRf++4lKFfhjKnaEsqusRn
Xf56RAVqiFZOMOE0sSjUE+wZMx03jm62S2wXHSRqo0tYBDnV+5yU4y/MO1y8/Kr1tgX8lvQMSgLj
NP7JDtxx8T9xDf5WUaTSkbPQr1d9vHYJvi8w09K2NiyDAJfcr6cTkj0rjj2nyVtwAAlKcDPMZaty
MGmz+AAQ2QP0xYiKQSdtdvQlxE0/wVdLax59F+KAHxQSl1Uwfup1E9VZY5c45NnwGdKZ7W5zkRgd
LvSs78WwKIkSmTBvnwP/T2m+xLi8MLQr6h6OCVIQzOwIz8BfDn9lgAE1gBLTL0T877frXt2aGcyF
6ocFWAGhmrkywDy5/4U/iXMKHix+1w0E5o/dPSP9LaqHDoJU32IikoNuldUxckw5/9XHdqUEXD6j
/SAfIL1aFzRE2I8zA4/jzyv0F1EN+YwhmZheKVPW0GScnuuLBiGcghKoLCe7tP2NTPA59vZEsEOu
BBL26UDD3A5Dgm4HlBL2GatEAbeo1jrmW9zexPrwdGq6DW/kVpNe2acbvXvj1g8rwFHbjo6u1TI5
Bw9zLegk3gzxC4EWB2WH5h4lxFgdezx84nWiGutydAeObZ3r1WqOiiCzVdcrYxyEeOHsq0tWoIVr
vpTpN2x+NW1OxEA5xNEUKfsGgczqAwhxY2tZCGk5+k/X8j1jGv/BAe/9x+b5mqpSjVrZAIWt9WaS
M1F/43w5FkjOsW2V1oXSE7mxoqJqGkdh71SGHUkGfUK+PY0lBx/iZ3wu+ic8uISjHlbrsF4mEQPU
xCGOalmefX9rQ3De+QV12QVvMC7gnZ/EBiz9fsjB9yf+x/3zBCwron642V/unDrPLOAF4hBOrhfS
2Bo8B7WzvX3RvMpgzgBEPVqlfGA92QDRjgcMNpOwZ4qXOFjiCjezZvt+MKU0GVdS8XW5tdNg9ray
awD7Uek0yHApZibR3RB1QbW29Ls6NSdJi1TmWmroxU/k3azn7vO+R6CKYSoA13OdcgSS82kH89Mr
ja+25JoKbgISwb2GmRWhDL6DXhKnU9tLI72yhw+lDVa4DQ42tPv31jahIvx3YAY2sRY6JuzDE3C/
ntsf4/kLPxj+2rgOXT8YwHQd4J2IfmVmdPlMRmHs8jqGnu+m5rKqL+MVdCeGHSA/05rYplIJDk2c
2DJuRE/ldHxUEi6BCWBleDjRSv6sPDxcex4mjMZfJFQQUMSkB+tM7uEHrCNhgWEwQP4JT3QtPBIZ
jic5UD2ws9Sp2DfSPUSXqjRasDOa0wVZu8v1Q02FPcCyWDgbxOhDmc0Lm/FzphceGhx+wzr/Q7eY
Ta/NnMyJ6noTwsiG1CuoGaqN3xPcA3azKkX4NUjxSBFHR5MqAPLeIH63A/8CO6gzKKp5X6gMEwem
nddFat32/8ZTXijjdChW1tqj3aZqJ+2y1/oIu0KiA9AgNkmBFAaaWDoJ6Z/E7e/vwJ4Vj3ajvJSR
uM3K6t+PXBbETWJM/WOoiz8L8J/YrOeTCHCircV7CKqNi5vhuqqGR9Vw8sNCcw+LykJwt+39U/Fx
sKjbsgtmR8X3FiaEdMqdQ/cr83Ql24BqEbE0izuI4qiOVwvViZDIgdOMWyb/RiJq2OxJJ8F3ZlK3
jQaO9qe5vKm5wWucwUnA+uCVO5d5o2D9CZFXCvbKTEXMCCK4WRFxN5W/AQTbFlpTO4BN5I95Gno/
zEZAP8XZKlMk+2XpT8LflzOYPeQqoqGqDAsN91+92IO8iaD5YhylQQIhLKxVH47h4vh3ydtVzJvD
RHiwAoaEGjq1Bv+1eCnndJLcOk751+4VEB0j+lM4ysUkZJm3HlqiATUq2Ta6XFOFuw98MZ83NBKd
Pxr+Uf/wLyE9offbvAj9uTS+JRvh8r60jSmGbE9fpxFnGL8jMbQeiaQn6D5EPEtP9NFNQCu5O+LG
oWpFxv5HOQkdqxxOZHU9nWw8UKW7MaHYzVZtgdBgrWY6YBrESjTzM4xVodqhEjf9HGJUWXgl9/ey
BJBI4M6+tO0L5V/RWUKR0gDa6ZYcBeKmA2H5ARLmx6ZEsSykHqTHHPGNPp2i4uVIzN9RSAYjekul
uum0QZA5sN8WUpjy6nklNyCh5RmLdB9Tsz+bZgcQevczbUmYf01bykwrtoMG/JSXzcjWZR+gmEp7
FqIOyB/J8Be62zAeTYtNtIeOg0GVYqqXm5agxHLs4cQN5uFoTqZzuF9PywSZ3DgAWGqfpXcjR1oJ
BfeYDUtW7Mdz6AIXJAwThIFLkXGgDTcGKd5bN9KKxQ9mUeDvagZId/khPvXlC/iuaoLe5dir97OD
LndVG5pojab23pwh4mKoCbfE5mxwTVeTTmcdU+MCEalsPxYZD3uduanMertwrEjitZYjBe43bLkx
RBQO64PGE5fmlaZ11JOsGQlmyCaImMOQvzyxYs1X6QqdDurV0hKFxtgfUa5oKIdhmWPi7eYIODcl
K5Ocmzjbjh0qM5ycaQSvgiSNQqa6kHw38TwvQMkrXuwwPTx1lVSUctSPXroOtEfr87ZDzqVovlCW
Ltv5OxpFMCpeFyNZDS+0juU1Sq4yyyM39omqMdPTPzsP5awlgXK3wzzI30eosBL75SCoSqf39nPS
2CL3SIcKUOUF2x9ixkGlW85qv0B0Ikkk/GbAlf7SLaBgZ0fn+s+rLikCn22dyRoGoYgaFB0yBz8L
rQp4/Wszllxjee9bd+7D8kKDCJv3a7KPavh5FwrWfdnQgokYYcfHQ3Eoa664pmPBBK9WcqNDLGFb
CRKK92yDpsAiEiACoSa/l0QfPXEbzCBIgXW7D6NZ19Vbz0yl1Ec8Xww77ju/atV9ywMuCcKDjUf0
z4rrogMlYmV5Uifrwrf1P/c7Kvb+hl24nAX2WvZjmtfjGKMR4/fH5IRRkHCxFodPWmikCU5Hs3Hm
eP6+KU9njkYnc/2fxqEzFfBdmuLb1fjO6VunilQxFq9jqwPWZHkgYSk2rbdgxqfZ8HpLSrxS+ktd
XOPawtpKYDcqRrK/OPqbGIu3NIMOsl5KXpzUCWxV+VeKm1egx8yLDh0nu+bSpeyfpR6tkT+fsctl
lHrqbT9i9cUPIacSMq4aWWIjWHQRz0VawtphAC/1RYUzYqgK1f6WwU7dW2l++OHav8SfrzAa1e6H
stdKHohUII7RkHahrGtk4xvYPdoJ7m8Y4cgNNkiVeNxH6f4CVwtblorz+wjW5FHqY5ACURQi/xEs
xlfpy5MUwUPqbeFilccpegnoHJ3c3qCV0IlkDE7HUGx7NiNiL30CVvU4kQQPUIrQeq7FL/fF+xqy
yukuNH19pvxANGtWRLWY/ViGO2jZr7osPbmCJnRuwMMdb0v2nKD9q3xBGQRa9CW4SyokekW0bPlz
DXjFVfJtz28jzEGXUnM8ja7kdoIWIG5eZTfaB3OcSPptZT/iI6XHsp+luluClfyvPiMeD+wxv2km
JE2un3NhIuBArKZ1wo2wJH97KeJJjxzkivoaT5vXD25GLkQ6rUUTbyaCJHiKNhrrcf6e4k9Wl5x/
nG3m1SIsVWoFhBk55oLuQ0K4G9E/BrKfsXgjs2fEcvNrj9A7dJb5zRayjo2IkaTus4y84dwEod49
ncFyAYNQpGZ3xRwACQlVUoxCST1w0f1aOBmJVvacBzVB8vgDxc8LuTUKvmumRY8M9GjPTNuY+syU
yG5h5o1ZhcNr9AEs2uDyksSWg1/mO3mQ/aAGss/+8xdmoSjgAhdFxPxBpM6zuKYxsmx5gUt/Yx0V
ChynJRjxlJjoiz3x/N/a8F2kjP8BK9onU4LqL+/1go/yp+mkPUIPs+NSfUXMC8E7xLuMA19pnRO/
m0usINqsb9kz6Qg+U9CSiBQ0sP25boYZ5d6dIAwaeGwzQrxR0EU8mpECm7L4fTQ2ydorSZmsuzmC
DLGt+4D6pA2XFO1ARmW3f8nundH5/5xwqRaGUvMimQE+Qx6P3+k1NE8UPg744r5y/XcimkSfFLUy
sZIeIOdOLFMXGl6hqltON0mdFED7+mdU+A+uD1wiXsFcru23uT84WEJxVURPk7wZeNfrs6EAmLVq
ENa7PFr2jh7DtjcHLXX75HAVJr/VpDLSDzQeuPCcvAB5w/E3txZEjAIgQwfRoFDyBszgat8Duxty
MsYRjsUbHXIpuOdPTIWN1JNsdHjV5WDDyfs4FP9d7/dmukLKm5JzzvEWfdtRWxwOzEBAZl6NntCV
xMfHCn0aE7URVO7LHfCHszMX2qaZJgRF6W68CP8txCofRqmXX/zj4uMUbjTmmS69V+NxCqdAV+lO
L8/QtB34fD+FZ0Yl8PqBMjKh8rLcPoG6RqI7gMyNSZ4IrxVGxSYIcF/B+hjnbkKw4tctdaKZs4uk
Iv3ZPi6CIpGpmAVFaAoLIjmXNkzcfH/hMFzLvE6x03HkKYovyWt0pw2ASg7JsH7kbk5YqID9ZGff
Cp/vIfqN3G0QEsXnMRgVlwCcRnrixHVRa9uJ9fPSyOB7awzSaulJ4fGZPgWPH9XUZet1O2ZTihV2
xtbLLmQowlfwDPynYQYixO+ldCbDHyES+fKMSpfr1EjKasHCs5KyCvCxrIlwWX5Vafh//1chSFLh
5CoHzHLo1p0PbuNHz4dV4hkFifqFDvkwNrUS8d+JQUipaYH33uXzeRz24tcfeQli67zUWRRJWUm+
qLAfJ5pxTe8QdKOR60hw5qQJl4HpxbiHGMdgs10041wny90LE098JX2KAvnguHt+9hPzYRy1B632
3BsdHphXRIaX3OXpI275M/j7OzpEWe+OXsCYznQmeIVEuAqMok6F5Hl7tqhBm8iJeQq/UWG22M8e
uOPOzhV1PKJgnqtsPrgkQaMr1flcwh3BmloZ+WvpnNAxeOBi+ruKJKsVqjOrrFUp3btmBG1hDQb5
m38qtmfZf5PNlV3vgqpKRw0EVOFI3NlBLeylIXf0vhMkgEyBJSDDsb4/AccBEHOwaFUzEcuPVfR8
rz3XyrtYjH2OPJvJXkgfmcdRWsFwrhIk1Xw2J6/waZszp/oQWa29iIQyvXDFWwjYrcAlMjhcuKNh
D+uWXdvyx6K9jk3TCMvyXOUFSZX7AZ2gU154oAq7wZQ80s3rITJCSJK/utEJ34GYjX8KAFVEx6ul
boXw3o0caVd79VOWDX7NI0ufQxwgxaXMtfg052oJ6QgNy9wVOcQB4g90lqy0E2ecwrcwcQpzNsL4
yqB2frP/RzF0mHJ27yV9fWmxtsm7YQswwPJMsT0+f4zIZN5JGeNBUqEJXBDHhNW546rghy+5neyy
HJdf2xuXoPjLZvJEucx/BJO+3n9eFfjHT2Ta5woid4+SiKe9CGUFFcPUmP0cAphL6OHPemz1edWr
oPf75MGZ3JftGQq4Zj4rWod2ecJeDqyb7IzCucZ5JPjegiSuKF3Ag0BG+/gDRs+Tl0w5vPIYbQmE
7P5iDxjt5rOyWiU46Hmb77IXfi//TwxWhAqCIi0kY0R0mbqZ2vI3mk+NczXqqhjbNLpnfmxxnLwy
nBNz/cTTFQ9GXhQN8d5lVsqFS4nva1PLufIf0+GC+o9yLeIymPI9YCwjNqsrVCmdV8baZcwsnM+0
/TIIc5XeUrNuM/Lux9khBDf6dMXAVAQgliKX2pmD6JPWt2GIyuCRxasi6QsIWXWCUB0uT6dtLqLw
hvMjEdb5D6odOLqt7jvTZWmx4usI0SQ7zIgW/okoacXGjkJlpfM8N9D1F439qzYDe9/fcb6tELpJ
eKO0n5LdtEHoxHt07Tfv5B8kfeM/eUd07ukdu1a20fEuzzqrwgj5vVX56ueZSiOTA0++5a4YlCP2
M58T/1fdTS8O0JzwoEPQF1yMaPZ+VeOvpY4LODCb55HEZS4bGJRR098UYLrGiGz9YY9DqHiK4wkm
vwQiGqyQVsQ/fZzWodR+O4no2QiH6dmkMHYhGbtjEpEF/lzBnCgtDBqZ6/nIrtzQJlcGNVFLtFkQ
eDraqiAvp3Q9+TuduDJ17KZ+oy02Dyr4RWwpXEX5qq2Ths5wb4894FJsIZrNMvtmNqQfkgOg8guf
YbDjkFjhhDr+xGM57isRcfvaXPrgFcVBB61VzuTXQgbEEDOQuTxOkMBmfE93lasYdEnqDAcw+yfz
RtatPhJEGYynzikmIyX3sLQzGPvwyX4TGkkMQuC2eG2mPuSnMkfnze/duakC/cM5yKYWHjmEO7Ns
RTCJJ+/Xvt6qaNHFsBDFv6pn0fonkmLxkUOk+qELefwuFl0emS+zhtL/JJ3jB/DN4toqOx0pu++Y
6Vt6l9Lu6UtsdqWnwpLfeQg7Z8Np0cdHwKI1SL8Wj5L3TC3NgiULObudFmk9ft/owh2dcrxkfkII
+Kqh1aSGAvsu9IFZHm4R+Ay3zFOQdv0Wm1WM7NgWAykz8gU2K4cHkJcqFqiap39vegLKMzgVvBcE
8oQGualAtUbSHHyyQeLcnmnPK/5Ag+a2ZJeI5Lgry09LjsR4V7cucJJzL6pcZQASEARXgstEWAL/
k8Q3tAWuR2WZNEGEYtPSkKywR6K9j84CmtaNYJoWAkgdTfbZH4vDYlm0E4UkU6PF50b3UGMG8Ph+
ibkgbZt3WVdVeGLTalZPUC0Zwi3rqbfxE01nFYrqXKpqcF+PHB5Qkr/RFSnc5ZpxBqWpdIq/xHw5
lid23a2MwPJXmHpDiLvdUl6ZDaBgRr/Rkz6V6f8da7K6fnUH9vWAmW7tuaZExpdxNAolrlXfPw9M
YwvuAsB2Ri22Fu10WKMc7ayhN/WMlSRTDas1A4bE/RfcVHN2R0D6ghkoDxNsayH3bpjQoRoik0ux
aU2dr5h0w7h7mGI+/i25ZNoRL+Uf6XoMjOGdwxHsBvAFD//yh7RdBhY5tRpA89pkFXTXC560NQyG
uDOI+Vn0Ka24nm52ZoMU1ffb4/bs+PaujjfnH0EXWOBHbRE5saNWitU/YQz8w5uR9JXHOdEoaRm+
irmUb3Ky5E6P2lPzAC9m6hkVFTEphgWzOtMNYvxaOFawNNOYavN5KMAeAO6zkg+1VH5Nbmm0dUYa
kK98+I23SiOwxdxweaA9qaoUdaYl0Vc5UeC6t4EcTSQd8fIwoJ8XDcSdaVShJjL+nRabfZzs7CPW
jX/tsqq25S3SJBwpxuhibk725o//wNmwTGXPGUh7A0dZOTffyD8iOPrxX2nAc/JcrFDn+/h2VsJ9
6I/m+xHiN0CQDmW0WmziuS5rkzbc+szLzanr6+RW9nMmragt3wj58HqgrFDjeeIX+JffnB2uYREr
aY3fh6+myKxD6qPMHSqbD2VVdu2y+9QgJ3SPti9Creks+paVqFyk8B3RZZtJgHJo7EOvOz3W5XVX
DNo5rpdNu38rQZMrPXwuo4XSkIlWz05oP5pL67H/OPMhc5S1knzwQhqPCCfspKTbttdKEck8M5Ul
kAh2l4UUb92GYcs+kfYDQKUaGcBq9jzHUJ+UYnogg3xOTt/5qpIMnOIZd/4t3q9zj7aAnIq3S8LS
eBXKx58F3qvB4Qdl6b8NpGzVRZGMYNGVOePO1RoD9fhcjdQijG2NA/0D/XADW5nSZRWm2DrhtMH9
G8XQ9Nt2LkPKacflsX4SJ2PKuqA+te+gnobuyJKU+hax49mTxbbeim9u2nI8ptbpNubaPZLsQVuR
+cw5i+sZSwUHEeo7fjArLZxmKHOBBz6oNbji2x6xqgR/vKejYFn3hR2Nn/2376n5SLGvUWv4fagR
l7QqgSIeCdlvns3SpJEgM0zrrbjjOsnN51st2XXC86EyxY0mNwX0DbY74SjbiTVY3rGcRfuTMXB2
og2CIl3rqFQ7fETmmbQo7b/Fz9TUHrnfcL3LiE0yRjn5kubNY5gLsPdOWuRMzAT1H8MoL41DQP1I
u6K7c8u/qf+ZV36YhJe10AlTUbM2VEFYqWjBYQLugr1wSgkAJTZVf2Slsm8NNsqsTGiMFm/1caWt
AwpKm3iiJvNraLHloHSGhffCqhkgltQpnksp6uALHjJW3Lb0kLONeMU7vOz3Q7Ah1LTrIFAZBx7k
FSw/nz6Qhp4ExHKvedLaFCKKeznDeG6uPAhyAmZ/EDENCFJEYUGfE0b+rbG1/aU9hRkY2iGMnFrT
L7xcvFHN68bE5NA71cm+o3nQpE/6kQW0LDSDhrEqSrMN+sLlW8ukWuKjXiY7M9EyMlRmfFwSOg3A
5/YkMtcgQC5KnxjHCkt6LtJggwTZEfCIBGdm7gKejrZwjs8G4pP/DDP6REWYXdWIpWu/fqeiHja8
K4BWDYpBN/J+DTWCk1Mse4qt2igvsVU3PFwjHFpHeRv++5roLGMdttS/OwhUke7NFEEL1d1byCz/
zXQpRm3es905beJG7aZIPAhNQ5u1uciP/b9il6x3sb7KE+cxoXF/n2nDC2VtWL8PLQToaZcMvkMM
X9xBzhgt6U4V6PmxAPYNEv3W5/tjtI1czl1KLQo8/srOdWL6+qp7HTPj6aREouVZDNBg2htuikRX
9hkfmilTHYqz5ld6hTUlAmAVF5tOQ4K5VNffmaFX59W4wncFxOpMh4L90fvzTu0/e1RryJhEhtZr
kNqiVO1DNLjeSdz8609sw4ZZD2vS1oJZjVm8pbpqn9PEO9pHPOrkF+LYsZ4DBtg/0A0eS0YTbwps
ky5ezCzeSrpjtY2Z/WKTGINyuMGB9s09EPXtIjtm5LmSIAFZbc4FOaHDr6MMQNztvAaHS0Ohsty4
+lkR0RTW74S5bNwyDW5ucKbNh507lMlfsixejCPndEwP/uf2psxBEJAD/E2qcQbKgDxZ9iz9Yzkx
uawhNNLWetQFDzk0dVZw+Hi6OeMWjy7Tuc8/TT0oFPiUVrB9lFhyHx0mVmf3ePPJqw986mxZ6ffi
QqGq8fCN1oLu0NeddaH9vaL9fhuQByEoMouqvKbtjmlaKtGNJL5xz2nTYTsEnnCHuC0oDU5C5Zaj
nJIwpoTbfAKE0htDu/Piu7bhwbpWojnkP3SkX3UjPhQuFsi6mH4oeUPvfsXgkeMfx4TB0anT4fb2
FcU6iocjlPFpTxxpJ1Y40yRKRMRTsE9TYai2w2LMcvdK5NCJz8yHASfwsm7LjszYqTpiUEtpZE++
m8nmWfIpiIfwVFISvjGm2YXaWFhKA2LmR3rIA3siknlq2mhvdylJWlZqI/MhmYuIConuTSRcDAKB
iCTLlj+wo/fLrbtBdUrM1+uUyCwH+xbmRYUUKLqr5QAYKck/kf1shELiy7V7SjGsMJFQI/t3W4A5
mFSM2u4SVrL5LDyARnlCmscYaSnf6c/SNGf0TZmt0wbaaFgapbshdt1aACPpFPs/bYcOJAiPu0bY
VjDOQQltKD2jSf9ZQtA2lsRyQREbSBNvrErBUvR7dJv6vxWXJoPAQI0PoLhPNCARdHG1nEpbHY94
LjhoRCTBzsUsHpZCmSzmw+yaHNYIvGdG5zzypP1mhIcc7YV3ohMx/KJLT5ste7xMa8oH3dKFQUHk
rwLplA9qSDEqjIXYu4HAY/3k9UPTTUtDgRymDpUH1IY13Ciwxv2dgY/0Oa6MGBwAkybdpfVmMymW
nna5pdPLBYbqWOgGbhM8JWrQ5SZ4TagNue3eJYLFwS+DHzOWTKNsfZLy0LaZQ9ke4Izn0kzhKSJT
HuT2Ttbg0TZxeB0lHMEdU5MwNLJLX6kiIKR9ZreZpRPUIg8OKA2gb0EeaDx0je0j2gVg544riMIZ
dlS1gRHUZSu90tmP6/8Zt0TYfHmTOjwHUPsAn27rAr+IWJnlIqi+q+KFN1UO9+3rFnPVU/vzqgsJ
dOIRWnrGW48KehExQWqppLCyiNkt61XJLLIx+y3Wt31DMQXpR3BEyXfayaem37Vbf2J4EIOZF1ug
rR1zZFGnxsTV3Q9Jag8HC+WzKk7sr4cI3ew42c5CBwkrpuWX0bY2unA/sjYFldAW4t8aYmHM8mLK
QHaOmZqzorlKpQ7oEB9UEyUjIklAj5KIXVwvnRyakwP1Pdb6mI48sLsqx4uUXtVa4bjirFjP3/9e
3N8mm3Ilt9VMmHdKgPTKrre467Pz+J42AsBySdxdmOsR9x2akIiMldob2GFuLOh0KSngHTu+cxT+
waOxozyqk3cTQziu9rqHkGCBJFwSx+02PdT+WFntC+fS56904N2pbwBCGBriUH4eHo9pFwz4DF58
Yhc/eVEyk28wKQ5KjunYApghewRlo7WnvhEAku8IUqqmgSJVb9csB/dQZv36xIkPmwZPpo6tbSHF
+5bvFUdd+QqmFDQv+uSQaSzgY2aQYDzT+s0eHy+P5vte+/5Jg0COsZrno9+tqYf/7GVznPYDGqdc
KKP5Hk24PIGcCj4KDKt+MrCNpped8Hs2D5hTBc/vQblsZjkbuj6O9NYD5GkJtlPzpnB0bhDj547d
r6sPa6Sfq+zjX2afkXOfH9k7HQI1QhpuZAjrfaSXokRdG4BkVn8zthRpJg7ns4qemeoQH6YgNhWE
9eSySb5YKvh7ip5K0Uin9J49G7oCb+TGtagB8U7LJjd1hCZdWX5dlQm6rKlCAsKg28/ZYgleJgW1
K3sxoxvKbGKGs+q+O9bRsn5ignmaFpVTaLxM/nGcdUP3rZ7n7JHfu15cvYT7bVo4d2mPDkZAe7Bb
e5sxo7JSVpSqoZCfx1yQ53bHTQxc8h1r+o/7ziHJLqvFV1TsXP+4Uw4kuxHhzyUplBR+kMDtQ4DC
QMU3nbxUFEV2BCuxbtC4xobHvMgZB2pppEc2mnTxSn2x5h4OOm6VBiy4ugh08Z1JaabwF8HxGV8U
ga5mC4/ewX0lDhKvLaNExgDyzqdRg7Ql85/a8yZlWjECWZ2kaXzRze16SwzFP8zO7q39qgwdPniE
udszyFfYR4lhPhpKeLSe4JtskEjqxwQsJqzhoi1XLZzzHZBKd7mMwCjtZRNlBQvoH3hsqmeItRbG
w/u4f1GIrNCCsMUfcLp28xIFcUI5yFZuJlVNtNKgeT5wJC32scHb3pmXjqIj+t2RirSAVz243+iA
w1x3cHuswTBzR/I/lcfJj7JPxC+FS0dhJut/QvjDvA91eHywHJEXowe15Ukhv7EtyFQPi/8Z3I2b
1SqkS6FxIj1TCgudbdKiActgtpFvvyIKQ5V1t9UySXpEJs0su8mhuFF/lSKyTzK2uuByIlRnhDcf
9LCcKvtHWdLjJY1RjnbmgFTrjJrimxu/MDg8feevSTNzsc+4WiIKoVfcyddVgF8lEv77KQvmLsGE
8RYHhy+EfPnEzGuk/2srpFjhJPP3MKySuI0FCRP4tR0OXwz5sEmBTec+q2lW1vvCI0buqSkrgE8X
K8s+vqDF+3bsfsGgQSeI8Z8GQbpYXjUphDMfOpKkT8edMqY0/LICqipefvVefPWeMZjgFD+nkyjw
4+cThJ7YZV11TG/8lVfd/qiKBTIw3v1vkYHoztrHIisFvnK6JTThgsDwLo8nKgTDwdtEDD5so+Ib
2Az4IzvdxKcohg3tf7qpkekjfPVV0H0FfhEc3tc+WBc8c+ywCsTouQ4ui8MCW2fG2V6t7eyMo99M
8rJkY1K8qLwQx19FGyAuOXoe97ZGrpgfeIAGFgafr0vf8idzAse9G+B5IX4nmDamtwxxA/4Tge09
wH66EkZhwCZR4QSSBSm5okhlCBoCWBe2xAWS5p7zuKRej2VFtdPLtGyAOdx8Q87why24HiCF/qZE
vR+2Jj2QQgIZ+ie13bgrCfaO3lkq8nDofzCmMhxRHCf2XASMfjYN8Co9E4KPz19XycgtqgJNlvlq
PbtX2/RKKfXSFGjlFH5zvfwoSE0Yzs5AWOc+vvyCcMgzfACluabSyvsXiCKjFYrWc3f8ARbcM9vA
mGQgR9CZ63RQQUXUUQjBst/sLVnW5YedLsVUg8pSBB3/kAuFypAAQlsNxd9+VodrUWt5aIjmIhC/
hK//AwqBYokT1pQQQIaAuiHfZoB6frowEfY0Nn/j9eGlpotBOKZ4fA42T7V0EfdvNMxeP0/5KlT5
Rx4BDK1TdHq3q3ZUNphFHSEWn+QX6iT48R4P3KDLYKY2ehPo99CSASihPsDYl3pbDX9bV/WgxiIe
IRbR6lgD+ddGsT0qHDfolR0F9p5BEZEos09oj42Yz+BXXR0CZjZovD9nUoD1yleNh7BDyAE2KkSc
97R+8p1KMkM6A7eDa6zCQtzsGAbaPn3Vbhhw1wwHJToi9WzIpSWWAnWbQP53sdQB5tbJ7pzY4ynm
XIz44ffBRfFjQND/3duFu3e2IrU+NoySeYfzUh7wo+ci2lI23iiv+zKSuwXbjTY/PKZsnW94ihO6
77UlSouIy9NuC+Ny8ZJ6FiI12/E0YeNlhQpeq7Hk2bQK0S94BYqp/ZHgYHz41q4KB7dpVZxy7kkk
DbDDg/+nBrlo4eUXIrpag6tnZMLDjUDmSO24cHGlwfT6YeVV3zytXt6Xtyth/jbh8Cz9CuJczgxU
qAeoRjXHGI6i7pXAs0b3+6E4+oMquzjr3mWnImBM/n8CTvXFtEfB/lEb38V6xdAgFVPOg7DqAGKb
9+a7vWZ1U/4hFP/4ym4n3ma4QQi4GvdhIXalP9ZeNZ1GfgieGf1Od5dP8lLXFNqS0o558E9RhhF+
RvsSv0YkeKetkK2WP+778o5yUw9iVrYlmZdZ4ZFdrzC58dNxDEwn2BmZ+GNZ47L9sax7cje+yHqB
O2nWMpfm3WMd0oVJHOy4Oo5Hz5Jm+e9iNfyqeauGmpmatHQg4nd/bFbxJATgeXgftGO3g5OoJ93O
/jLEwvq+VyBptKQMlFZz8Zm8C9ED/1dL99tpNOhPdfY2IbHj57LCYXC7OjqzrxZIUSYS/+TmKuYU
ToUe1NMzLI/v6xRJduzHBNAqJ2VEBW0XE5juiAzAGJ4vC4OsD7m/THH8V4jKr+0iDzv/UeT9DENK
VFaKrZ15FApM+K2okQrWVGrP1YgA0VOwGtxRTboJFox0x9AXjlHjRgF8hLWrVgJCOpbc2xRqpRDj
qpFlGxZKZzU7smZSYk9l53IWSOovU0IcAH6e16F1u8Sgw78UcCO1si+Wc8KKvd0E1Pw7qNWmZk6X
bFz7Khvn/PvYr4i2HmiduqR763UMo5ibSh09YuephWlpXcpaen1sbjHuP00PTSBqbkRHx/9+fB4E
MOZgQ+ZVwcD78/iJfUxs400P8SkMxCVdgcztzWwwCmJYcDgmC2Pt8W5Nxh/5pljE5qOGfTQPndad
mQcG/AGHUs0HZQrZWJIZtYSNce4Dfy8SWOJYqNoefsBeZgjfnUPhHvTrLhDLHZFHfY/K7JzAOkIv
4bNQGtGPdIvsbtj5MzyfyxrcazTYYjo8/0CWbhAafp8EFtadCc/Ti5KTj+VkI7KP7+Z5WKLzbcTt
5kufzspbBGH3ZuNJejVJZ5Wks+u6PnhvuyblSQyq6sC3YSwGSaYOhpnxefFQPbl8VZ4Yesi0Oeem
Kwznyi6e+xTaHsnBTSu2no4MI3pc/EAVGFQHSdL8V+BVsQGw/LbPUm3Itsf9cx8ooI8cIMEyzSW1
gVjzAZgclmAGGuatSSne7+Lej8oQBm4tJdpwqoYmJFMFm6CwHQu8Gsh2EOK2JgOr2A7CLAjCR3Sd
sueBLLETgVOV2w42UfmNUrGjTpjg4LDu+7W5nDA8QUhjrn6zZce1DQ2wvtoeReyskZa1Gqh9siuG
6+PR1SKa1hhezXLYA4UpKVPW1v/IVst0zDGp2CijlSCWjqAzvR4+7wGFRO+jFujrKJubWh4rK24q
5HF5I6gMq9YHn2J+a9ZfRb566tIhNuu2EO1vgP566jh9VCiLyKilG2cZ4WzI6rDAlZEXonDA/D6i
GRlm+SgVBKsYWbvHK83V8H85NTY7KjqXJvbW/lt+sBFIT+5T+q/V1L12wnKHzJpzBY11xvUV3lML
u/g12J9+KAUKH3gymay9n6Fk6H7pBacb4nu4gs3OtxDyqsN14gtg5O2xAlqZ/dAGeR4hLlpL+i4O
BOjqJR8tsqvkcW90uKcFNix1x8BnfpyXeWAfERXNkLKyBslXuPiTK+Co8X4Zqej26BRTCR/3UgO+
w6qNBuOSdJhbRiZ0xyK9DOoAYnq1mKn5LY+cTpBY0mUCkAuwSEfAiHsC9zuxiWeCxSQv5yawZltn
UK7iKiUmpcCWu3uqjzjKQKe/Kj7OX9vb1zqlQKE1Emjht8YEp1PPIArmVFqljVH9XBl8neWfn8sG
JiNZGfVoSNlEVNiSBthLbGV+qmCfu6FH4lenCZJfaTaia6WqdmaPHNSapQ/mhtkezgYrztvlCxVE
5L/Rl4f1550DYJ6HhxUqkM+wUcAMXE0b80JiEWqtd/qJI4n3kIelWRFfsJkqnJbhv2foPTtB1Cq+
VyFFkQwm2jCo6Pg6xuIg5vggsnLjR9PjajYsle0SJo/E+k0msZh0gSbRqLBJldTbBC89ZQtHPEzx
9PBJLlrk8atnwko65AjeEeE6urIJwbF21tl8L7zVoMDiaDABFZ5ZXOyGavH6qNIgxx1gPH70ePOB
6QaQMxavBb8nN7gBM1aZZfDy3wT8cRq60qhqAuZpIAID25GBtnN12brit9IXazhixjNGEKzgb6Ci
Onnmmdkh9f0TCRZRM5GbIcnGrDTXNfzvgoJPWFNYP0+CQBF1gcz3JJa97R7A+2KVJn8ghoRHkRYP
SdZqEWhgn6xD4irAaAGT/gnLK86tZ2c2pTrbYff1u+YLJMFj9kxrG6xExyFYvrtecvYUUSutnOgT
6xqHStilts9Bgt16zaVmcpJ15ajkypBPc5CZhFNkX/O+I5HtfyRVn+C9Ho4Brx/chHjaCfpeM7Lg
Lv8MEWRDqL+yVvvd6I5Rip5RAp6YJwsc/Zwc3v/E9EUCx/mbFSVtewrWg+YTgGqpDxRX9yGk5Jo1
o572cik5Fe3mk3mjijnj16jWpoA7bPFWYuGWqWtuvOqjgUbtOHp34mNT/n+7V3lFUK75Khei28Ae
WApa52wyVCf4BHPkGpyBMvf4qpIrNVwLVJImd/MZEGL9+77IF6jjzAhEYiSqWVTLSylFoeQXIB/4
RHLnyE11FbBFWMVw0/MbDturTF9bLwELZYw+Fs/tFVEy0PSmgzDF74W1ZVSRl20Xdsebb4MpCWTp
nZpBDjUDBbETugKILVCI1yqjGPNAMeSVvNTEMFlz19cERvGJwIILL9UEwlMK3kAV5elwVVGnhEq+
e7aBYP9knz4BaI9W1CZtbhMxxrQfMYcq1KBIcnTwGe0q6hfrmJPxSx5x+2bahsqk3oXBVFP4ZJag
IrnZaFiBg7LchA1hRRlevEMwHUBKxlTbylT69frjnxXoxxjuD2/1Cl9R3pXeEYooGLG8ga5xQK0J
w4OUyWrZSUI0BvvvhaX6revAxHrdPet4wmz3J7b4UzpdbeUxhmlaatl3VP95ewumTECUC+ih5oKP
Ia0Anb5AT3R1pirYYUVAmD/mJwZjHQQz9rkOQpv/rXpX4v/r66C+higet+9m2Ep08OmnHHAJaJUM
FGSBL3mRjM/Z9zo+9dkXgCmpndKHfZzg9pIWSeDkOe3EtmmMAaiigohLBwpnGACcorNy75f5lc7r
3qTo9nHkcOnXz9eYmKTOs7bm3qxSFr0vSr4OnLL3GOEw2xKvW9dtKNqzTpsWFKVliGTjKvMN+WKH
kp5QuPy+iLyHtE/65yui6SKmprpOlLflYEvBCrzW1MIRBy9Ms4T27/nQhGt9TFQFs2kLJ/791k/c
9sZYw3Eh/QlkX8JyT5thM8HyhI1vpcvuPVZswIp4VnRRTCF3/ygC/dLhiIJBzomPbfPz9pQJhyad
vFOBgPemOFpio6OxKrOkIoGGSlNx3bj5WCCvY95YFbvqb6yPxDTMQb8KAyiSpxn/z2XAei6HNkED
tnZ5iPUWUhBFFfEgjcwupKz5iZL+8tTV9qw9H7m3z7ROSfTuYu17i785J62PMEp6gyeqmCAakaON
INTC5KwZzJZPDxNts5KrEKjd19+WE22lOiH90vX7XIDW0vbe2R+O0mktz5IMwfOLgmlAA4Jm21dd
PwxoOANXFBUzbVlICbAHTNmdRpRrSid/WTBdMu94nb7mqZQGcUqgDmXWFy4zfNr/BGhHll2/wxlL
tHbSY+ov82dyj5K9HJPCmQtsKkktVVfokZO8POzYLqcNLLkmkD9F1iSpIX6ggcphau2dU9Hmw7dx
gVuPXcIkgRE9RtDmv2zzQVCX0bnEFx1bR+f9AfBT7Gh/9ZkEMzglkFIrtOJjvmIZwc3jEbrmsZp4
Bdda9tKlrsgZM0eqOTkLsuO9NRdDOQKVV0965hKokpnU3BOw28z+j8qTFXfztHFdIFaqQDTbLztQ
726Au/qPbtSiqfH3ST027I7+NZGYHkG++AUqn8raFPwutRZCtFpEX8oReMJ5tK2NBU9DEJsJbVm0
3wVwsRSfdw1ODhNkuGaTP/ITRuS0SJlAdwEmu2yhvJyIkeDtnXPRaL+Lpo9mKNqj/LYgOIk1ZdVi
Rv48gn0TdxNWdJGT7ZTfT418z7eCqLhwoZPMYx6bIYqEEuWC+y+CAQ5EJ+zxz6Qy1ToPFpzUr5xq
KrcQD6zo/i/palJZBMypcjAK2SV3B+Oo5uAOWn8SXX4QyyeJnLbY/xCIdPSnqEWSO7P1ZrvSV8b9
hExWlCY5+7RtyNh7BraF19vNziGtf8GyOUGRoIr/4mYv9XDldZLKDP00aiR4y/IhQXxEnId+u4CT
FMfYnBTeL+SNYtuW6Bg/5ZIN3KaKC8eNzyeooAkMHZm95LPtERu8zuv8de+V8npkDZ1bkJM4ay2H
7rdcUpfs8hiCqr67k0097sBp2dXiZXTUYMosqvrkP2UpcEKQq8jct+Bq8RoScdMzxAaITLTwXNOg
PoUAO3ObQbatEXx+9dsEuuna7yiW/fOkW16VrWI7AL7QcKHkoQgDfxifP3XyEU8suwyVRdhFJ16a
ZqmZJ8BCRTT3zjbLXfGcU8R75xzaHXgTEuTJVPHvibOE5QgP4cvE2FPUTLhiTG7DR8oLFTlqhTcA
xkrX57vfLB8iA1YvPl/70PwMbUfR5cFaOb9vTvhlXx/S+nZqx9BV4fZrJx4OyuZsNj2XKBBO655j
zstQZMj+agNCz7vCeK9m6mujPGR6I8waqKMX4b+63QUU50ZxPSJxRvDdfK/ixO3G5dq/L++g8WqJ
jzDyRH3mYtRoJwGsqDFFIwPDC1NL0e8UJ9v8ywiG1/mP49QNx6jhP4WisurrzY2d31OELE9CmG9P
QJtC+QN0kF9816zoAHwHUr7ni+Ww6Xx8C4TQjlmSwpYEYPJwU/lZmZD18+mAAAVhNxHbbFw1OQ97
WIoKtVdWbd3+KDowHK6zQ0ZeEFho12sWs/jwlIqUa8iUkkpcQxJsTRc1uCe+rVuRKb0aUZ4uReCH
ZxM4XyWGwB0Dz3W1nzTXnhOfD+Y62wObhL5Y1CNFAf67upPqtpF3zmCTIBdByJLvBzhZ/EqG8fwG
Xg5MeNIEI7emyNSzYIh7MGxPG2iowRA+MZuYfMdDNAL7KQkiZWCJucOZk5tE6pkdH1WkH40aOobo
tvTPii0a8pFb47uueuDru4/YCVPDvD6e1qf6DDzrDoCjtMAjNdp/wk3l1bErTn0R+QSUCkuLuC5u
YCYnfXQwqxX0ZXjD9LtlXoWI8QvnK2tjtvSNHbTN7XxYwqk62OKLkXcyuhN7u6UBUyWNOSFvU7hW
NzBH+2atfA6fNhQy8RTw0pP+Pvz8Pz1nqC9X5Y03gCPXofCdXERWFIybB70cPUMVHUbBID9du3mw
CXIhaFO+4HrVHCCn71q7s6Li+60SWzoTsggjZ3Hj2eCBy6JGDZC93r8SQuGjBBXiwWYkI3hp5xhV
FiuT7oDQETsfagL0NGXkfA5RWTtdzhlCtvgI+flRKdJgl3/hSkJ9MsP+X5tujMcSJ3OicQZtw03X
p953/U2AeohORMqWGYcaM4fdKe6kI3dpnKPU/WLnMyi4pRpD876cdfuAjXTniGNzra/Qk+umdYpl
D9NO5ijis3IcQ788PpPSG23EtEvHMr92WH5vVHgLoW5ZZf4JMFXnM9MVtSjuNYhURIQaJLsBNk4f
4NhYPqLSQmbTIdPh1icGdwx3zcrWe3ZmW57z5/uMgR7oCnkQQ/kHyjuCX33Q1/R7CSUmoCjks8aY
IHxU8LaKKWittsAzWqnUOhSYuRtuvN4NPStZgjlPukm6RuObAzARKod5k/VcVECLxMuEIFO+43LD
uPloeMz2opMZbbrXANXSv28gXvjnJY+jk6Px1pBwuZjoZ6ziERf3qCyVQFb9T5mYkBjtI6N01cef
mUJ0ac9trmXc6muak8EOXNetzaqiYFfw/52IKI4p4l4unEnHgYAzegVV+mGb8hxlyxp+WutAZD8c
GaEaVZMQsB4ZTcomQkfQNOT5ruiroHDvgn1itnYPmWfxO5rsp5bQ39C1m8W75ubFzVx9OiJ4q/ZJ
GOy9fx5CJTGOaQPEA63wUuCW1nJ61ZLtH7ERr4BvgPC8bfeIRcqJaungTiHz3Wk/aZ8zVfGasHiv
ogKT8k8aAnKjasmSV6nBNhqEDVftJJAknUUOheaqNHLg2VjS8NtoKXQUB/wRSrEE70r0Cd95xEr+
fHqu5JNZGdNmFzKcV5VVIIzisEEBcRZ6QVE+vc59aSCGMft/FAvYHd21ZQWKRDJN+OGX4Db+OlCh
p+8f3zq7hHoWWGODm2cNeBqwy0xqJXc3AP7p1eDQ0JyTmTlItMGHh+r85OhljNTyeSkcIRWY8zw+
p7NeDTB+ec9beAp3mwiMfskDUQfs4zMAJv/Y6sCjgCn1PKiPQZzBsBf9/HbO36hDec2stfm/PMn/
oCZwDJBjser3gs0ssYqqzHACWnl6AdwBaP8U7x5tWyMLQkFhwhnVawHbiNu5tg6bcgH4pK/Uu6GW
39flVNrNVKG54Ly27IydsoT6DJFhLZSJrrqBeQl3XwBHR2upBuILqpCvMP+HYivoz6MTS/NALvz6
AisOzjh+ES0465r4rugKBiM3TF+EAIyAXWxYkAkyzMIBbOdtk/CWH3sKdTr5rw/H8b34H+Pws2+z
is4zO8lIy+DCwiXFjhoI3DEJiUN0Rs86vftb05d+cyQ2JfmFjghsIJFLocXux6LW1VZ4KUbMXVCA
0Nyg+ZJHbdUf2st7XWzuAO1C3JyP8YPCW99LUVPPMbWLLoAOkKpNDxExtX/HsBSKfR+vOAtSOq2D
v/PRCnxO6cZMGwVVO7FLRvRZWhPkUsF3jWAaRJPW7lfc19hwkkDA+foDNKbS1Q4OpKnJI5tUN03n
pBPvo49yqq5IMcTS+k1BaswFZaIpS2pc3pD2iJD3vH9zZ/LUiFhyKG13B1uW4Br4NaxUwKMou+60
kbP+162I6YWH/BAKaTvd0ixULffgR/pdeq3xi1qXv40OMN1VnRmjtgxUVnbO6s3ftggNWF3FXBH1
vuba2083t73b3zLVIRvBg2K3k3IXQq1m1tJHw1ESBcSogQvr1aHOFCROQM15BP0HMlO30++uQ6Pw
9MdHLtfdt3ZrU0CH9tRNEQgC1CitdYYhNFiAzQBPAtTbWdUpSVSgPEljZ0ywyc/enClV32U48PP2
tVI6YhcKlKvXVCuUJrBm9k8iUpWkBylYeCq7cfV/RZEo5v5OJUriSl9/XccJdr9KO5qQs8pM+Ub7
UTWAnoaV6zORr8yrd8u3XWwh14FZTIS6sVQv6+XDyPdFj7AcX65IjVP3fDYbWxciaKefcdaya4lA
aX0G0w6KjJ/DUHL5xie9n2F1KwUt+Ns21YRkeUcnd0Es3zyrM6EAvYV/MBTtO6PngQYfXDZFJout
g0mylN0OHsDpU0yMGnN5pC9jEMyeDBcfvET86aXCl3pXZzbjSba0urdnAZYFKTfD5M33bekTY7Il
iOOukh9IVqt1Tfj68VMfaZW68aCuWiwkX3u+LNnz84Fsh6W4Z7ePnaWS4oZ+yNHQ4zDGK89pi+ln
2sWU8GcwKrzkTq0TlQyyl2dPhv8hv7fj8+/Wnh/WZfIhDlftb1h7JxwgcRsQ1MRChoAeRWgKsVet
+fAxBC3aiPDFtuAuFAx8oRHll1LmFlpnBDjrqv8zJIlGvV5/jcJe0hpnCZwqTrSSf0aa1TyaxPoq
E6SZCyzCwhejD7YPdfWPtKRURsPm5wZm0Q7qHSG2AKRPxpCCFAtV1DiCgElD/RJl+PZBLTinNmMf
KLC9PfhNcT0UeA+ltdiBxq8rzNlnXIPhqJeKGrzBQscUKXNR/NHTGkhenKmuQjPdm0Oxea9e4GaA
j7TSBe53MIIIsNGf+islFfuMadTnEsyQHKcd+6CLvi2PhYx0+6KHt2Z4ZUj55GNcw2/VyhtIREWe
10KlXklH7a85ZkKzhPr4h5tRj+easCwwMfCShHXuYfnum2nivxSvLU8hF9/k82uUM14a3DT3Ju4B
5BsqGog1NqHGeBBn9UP6FulO4JOytKP0JYgxbXEdNIiIw3/XimFY21dTC2FAQenYajiA7PGLnT6X
B5K9AqN4Nnb1pVEU/j8S0UHdC9GIe2aZeBj6znoH4Z1LHvZTYemji71xQgyul8u0EIyZasmuSJpF
npQcf43E5i6WWzdOBnyOfHicTRF9tzt+7210FJq5QqHFgWYQMRb69epLErRTOSYtNskE1+GCDlxW
leMn0y3VNOZTL7DqoER+xiWPjCXuj6gFTJ9dWkRA5whHdlkLOgOWjTKLDX2c9z3vTM6Erp7VVwSm
iKQvR+svtkZ2rLx0L1IIrfGsynxEV929TVFImYezRkHwJRxuYpjlMYF7h0hbsxSTHt3TY0jxBEFE
OcXOMdOv/EZFTWpB7yOzi1tyBpmM2Hcl2dE/SqductAGLPc6KJSBCPh3UXGy/vVk9qpz92IZ24Kf
lDaXxsFDmsKtLaw053nZtP3NiVsF8mbxArlFvGaIMPlhMea8TyQtZPDivRfzYtIH83DLX9xlIP+P
NqJyYNCxJIiZSjp3fQD9rb9tuE4x2jGeAuvmWXNqjpnjoyKagYw8UwhO1kLp0Mvs7VhhsDOr4vhd
NzyMRXw4CEeU7K25gr6uLPr9KRaLlCtcNhZ2DJPn8bgSqNSV1oE8Q6mUGXHhSPrHuS1Dfz66mYxM
7NJHPrqEdJevxY/4xqjwHambCBejGUz3ulgY17YQnCJ4d6PyZPVSKdZNhQY/EmXlDraZBFmji/af
+zoQgiD36i/ctoivJAr7RPEGqMjGUGdLayuXSDpZRyr8QWHnkZfJWQsNa36WnTt3HMNrqjAsBaRr
1qqF1WMYmRnvYwM7RNoFmT/Rjycu0HhNv5xNl+PR4dXx/APWTW2FwfHajpv7fMcmhZB6DDaD3NIc
pbHIaxgMQYtaAxpVxmpiPtPidkl84XrofuJm6w1Nh5peI5WHEB4/WTdInU/h8bjH/629WCu2xd42
KguCIU5I74bnQlv0E1ZRvtx85oMKnUnPb86teRyLktTKgTvd1VeU29gDL66W8w8dccN8kDh34x24
oDn+pdd9/tZCVKwkFfDKd7YG6w89CO/CB7+wsVrXG2WXI2akwNzZtQVw6xBC6b4/jT9YTd+VpYWA
lZzx0ob1ENXIf139LVE3prMpTtbczS8mDe0sVd0KPdmKHJeYgd5qXhWTdaZfygb+xDHX5l6gUut5
nIhnQfhbmsGPr2bGk0McXKZ7FU0uFILQ+ys21bTGVKn7ReVljfhKINbyI8OE0D1Eo7yluBbrt4Ic
RHhm3u7I+DO01F5WmuIBnfY2mE6rwWoACVcxDSix7CT940kDXvkSUXV1feWYY40umven8z4EzK7Z
2lXtAa8jX1ax322bD4tWw9+aPdSDWmWOCKHbxegnMbECcis9hdoOQHDan55rGvGFEHMm9NfiN7Tr
ktimRg9GI84XXt7FSNEZXB7EeWSTZmFkAqCw4TK1V2Ek1btn+sxa+CgEJxRASexy1EDVr/ajh892
lx2QI9g3uADCu3j68mMECdKKYxh1ttFMmRzJmj0qR4R2C/ikm0jGMG/PH1Fvkm7mbKv7To/JdLV7
w0NWswZtDAVjD1ddqDDrMEEY3gnlXFwKIexnYslC0KZCZ7WOUj8CRjWzUupdLT+ZLy11xz70RY4J
dUeeIQxxB6hRLWOOxuhx8ss4gqdr4wNvyiYaeCtKjdzaVrsMcIyxq6tp0jzgkxtO+NU6OD5Ta8Wk
dLTf77NUVf/uQnlNWqr/LKuZpvu10i4ObwgfcywH4FcUhaL75vVVHqZBaZFBQPh8j2rr67jlsN+R
zQOqq8LqpL6cXbxAQj7tiexZ6kyMZZU1n/wdhOH2w6K5KxqUMQ6X8SpG9YRFd4zWr1oA1Td8P8vE
rL+nfjdZzi70hhaBnEciwm6vnN8DcXEb+hjFwo84fdGpqE7uFbd+CuE0c0DwplMVvxjye1eWtyzS
lX65IYXDb6EhZU09kRo/fqXPlojpK5MZkn+9yIJp7lykMEZ+mYfSyslGpYLolO7ARVEbmy5vV3eV
5NsYevDmn7CUeyW4X+PBHgvFvv20ZLJhe/bx8tr5he5xhvDODGKo+36xJawMPK13xuxwsoQiutWz
sbEDQFBtzr8HSad7cRqwOrfSu38BlvuJY6QRsf14YjJWraRKfoeLvPSp2pWDhr5iEYj/uJaRrhN4
Ak+Z/903moDYG3X0tLPXZ/HoUoVnROt9SVwV1G05he1UTkl4n/G2C0exjvYxgDun/ts4KKkiFFuR
QSKzOPLX2v15En/gfrLpNq1IjfK2tCAdIA2739svT5PBjljcBe9GYAZeKXqcJn2iKM27qxezwahB
b4o5Tk8f52/U/kEpmyWo/10+eRN6wfSo1/ZlBTy3x8sh3rN7iAI3Qqn4MuoJYjCyFlWxy656ySMj
eM+AFH74S4CjgxT1mCz37QN6XVCBZP8OoL0DTjb3X3AkMqk2jfMj6zebo+W9k1GweuuNTYbiK+L+
lLj0Ng4SWsRy0BOFHAxRKdGs8OpDplSBoHiaJMNeIaLp58luwTQlTiMyWhJeTQY1AWTJHlbjFskv
k1EN2dx9JYjRz8gg6k2kHNB/E0BqGqOpyyTPj6aw5azcE/S616CcUE4JvsnWdIq7ZBvHzUgWwOXb
Q2ZAaLqaIdnwGX1hQv62Z4RML2ObEny16wVfrOcDqTb28RkggByutaP8dvPB2oIJlaxXQ/VL/98O
56aHvbvIU7Ogbqjdi8r2v1c9riY9sDqTNivjxROYt7+Hi4EXO0pqn/vLjKUMmCbglMjb9hp1vLZb
bd0uWF2/zosaJj6OK3Vc0UsGYNPIWHlOxTxZElEAZH82WAO8wcasJ+3O4a7g7IcRHjP+Ur3RFq1h
gKipYfPE2tMEaFx7/90SNXeYTn3HkXcXAIyn25W/u5mp+KM75z1/xzfcfkXiBJCTb667gE/AenMc
Shj4kAY4no6mVIhbnHwGXn+5Ia2/0Bpw6+NFpQJf7MkD7BODwXkNL2n31M0tEjFSYbMEhc+ylNFc
aT6iT3Dv5or61QGJW9uhrOXwPZwePG9+aGpCdOqPFmhBhpdEUci42IlrF29eeLbAeGU2K5q7vXuf
WBH5SMt/AI4ygceUtQhh6rw5bAwJaMOm0iZ2Ii4bX/Wbsyk85hm+ZyTfqwzZaCNmdf3/BjyNG2Y9
K6yfcfSxvwVmlo6DjunV+50kMj/jFpeKg96aavWXTXXRL4FlNqdREKMBEC6pmpvhySIiSCGkCccH
cS+3/om9xJaqd7xXXjEMP2zwlTS3sxiN9+Grjykd+nsWh6yEl0GXlnramSW1MjVzLaYFJIaVZ70U
J2dmqM2mSSjGuHHNUalbO2DxvvHk2EYYeratlJbPGV9GkViSr6WrOPl+91Zgssgi9uEgYZx0OGp9
oTgjEVlNwUXrluyUlV7LUgDd+pTKZa0t2n9BfVrTIq13l5Xe878U1ch3IdUKbT0Apw1I4ddBs/Vo
mQgE0uu9sRIScTb8fqKMFHlj2pCjjaGR/DdQyRzo1xrzy0rN8Boh4lV0aciU3qU/kkJjL6GC0xDI
gB9QjKjhIfvYY1lRnXiFQGXX8L2tFKS2JPNZLSRBJ41u/RoUpHZ+SdQ0POoRK3HZDq7IWCh1kR8h
3PYMsvKT73DI6b7Sqbzzub28A1h8aE4v5I8ZAQlb4fyMQ5LMM8+iGsDi3vIej67xq2LM1Kj5N3bA
kG1eCxU1nfdDdqKbEmNp0jP7hjlS3pMhvXbZRDYPr2il5dGJUyavu9I0AF2hTuReqVnBVjcd3hF0
hAO4k94/d/WOUZUA8dXJprKsVRxxz6VylJzwJwDG4rBb2sxDh3H6DcElQ6zJiieI4C7LyGxfm8zB
qKeJSK4na6YziTXk+j6R0OlvaNRT87Z2G4He/nlC0k+vnMLtX9c3TPbK/t9i3Irvi98vG1zbajWk
lDXfUq8CiEF0sIkvRRcTfVgDh56/nsvRd2o4/6iYaNfyjFuuSlQ9Fspodbu/SM7+G+DLYH0KyYKx
daULqcHQYSfvWyImN/vIMeKmziQ5lv46IJ8c+ZMGii3VBIl4+4CE9uxMKDK5HhsueLxynjxMXC/0
abWffpJBV3hcKKPf0F88yRsltk/eV4UIRw8VDv2c02SGGndaxLyISNFxOMArhx+hSaALIDTHz3TA
FfmsWo5PsvWNzJn22bp7I6Sk5YztJYUwzJNLkqdOi3TLXIZaTpO7KmHvCdcIQ5kTCcCS0JhwjkHq
QrJD49lJhLhlLFDRc8X/1ug58McAPjX4j6b58VzgWLzv4NyyHr2t8ECDW1O2MKfSS6wXuIOQlkyN
F1GDfxAUoMQsn0DmFV9tkvjb2bEEkw0gLCwJbfIrHqJ4CD8pO2kPUOUvA8GgQlCyHLGbLFu3jCR5
aBJR5aMHbMwuWGpTc0fPOD3jqvaD23lVvUqQnp0HVpvnAytC2Pxp4wK5/DibGcsBdMVqyWBBWi+U
UU3uFujKWeT4Q8+FEaQ7P8DVnjOAYvvX+GIqzymlY5L/lH8G82E8VCype860CUucs2BVdsxTk1V+
DkkpnhF5SRRtBEIQc7QRuskS6O4Wj94w4ze6MPAwe9qONvWIcyXQ2vw6Y0tYw+xipquchsPHZFYX
5+xe1E9vMHEGufZblZpjZxN2MNylfzXDBXf06yHSN2TLTUhZEZjFCrJvJFJmFaWjPHlGXE7eLOGF
RK29I40+szFfIni8JjrqvQXmziKheDMbeLth2VXaCNa3+mrFdwq74JMQb6qUxA6PiIsb/uTgEBqn
YXN2F7IBW/rCiMq4cojt476kmUP9jlYffI7PYg9ot/gX+mebhh1D3DrGDSE82lqs5iH9QZmO6c1o
ybv4vpDOUgoh/2GH+wVHFiCAtmlBXKmyCVFeiB1g8xCqt+MTsQWPIhBJpWDXl6taEZiqrdxzfMyJ
wTx3wnDz4guQeVrKee/8Cm00vlTkgTex1QJKl7Ieox2H/uFSmY3p7izYqi6PlZSLDyr6RH209L9z
xLwDNaKbi4Qh/e3fK0a9uIpYr6yghAhUws8NqGdOKJ5eJwXTCSZ/SQGm1qdz4Ld/TbZvuq8W3kBb
vKDfeNtwHDzQta4NksUtiblTWcmGSKuzJkTXHKZEJO2X9qxfLByNQSMR8mFFf9gV0nzrBQob2eT0
rtmnY1jdXUcGi70QCojYbTmOyVWEJ4SzTcN9wN0ah4gCwMclxIhjBt2PFCJu7zU8zjk1pFm/o4N0
ATAPGADCUnlynZ4Py1vr1hU0z/nelB1uBxPqotFhPqPPOqnztvQDEdBPKRQPisVg1ZbQ4a8WRww2
x1oYPw0xPqi3wZVbe2kv54n3DSVUNAM2q4S0OATIc6MHdlebAs5kgcfwoSdxNsZ+XFBRzUy69TEh
rqurCD5v0YELIUsDa2cqKRLrmVBkckP+R+pSDCrfv5Vjn+MHyVfikZusLa9jorSZQQvy+PcrcVPf
ZrcZLaUSa4Ja3nMbP432v+hL+CSpPpTmpHgZdcUxrkIQpQ5mC84pu7LUTlpC3mcLxsfHvwYUxzbK
gDbKlWRThI9NR5BcOafUOcqLKdRyzmxaUth006KrVMiHtz4Rxhed+bJ02zuKMK6sdTZ6GKAHTpqI
s4dXP28VT9yNehZwHUFsS8I5ptNQh/7lYWgc3n6YbBff6Nk0r2JiPGQQn8VdmIub6l7TaPr1/HnO
xRP9Ko76TUq8JzEi6HrNZ2SRyeC484Ngc5nb51Fi6FqS6dvcJS0O+Cacv0T3oJQ+D36TSsIn1Ahc
DZovhQ8enjoxqEV7nEGeLgPP+X5JSeSgxbDMkfozAh2bSzfEJVh+R1JJp4n5jxr5Ul375CSFjRhq
HXwQWycKOpBRYuOvhgpwxMToL744kv3yVaDQ99vdyVfWrD5YmDTnWv980tj2mOOEMd/mkB8ldvTR
0Mil7F/DM2BNejys1CslblwBn+9z598SjQfVOOKSsYh3oipGiVJL0wemOMyX3q+bnu7kktaucRrw
/Ug0+HvPc25+iPd37Y1sFnoxj56wqxrBWhLgSnnOrIUnmZ3fIh4Kz/6IG3rXCGTggTmohTfo++cG
//z1c560mBEe3DW3QIO/eG/kKMOHfG7YwD0q8/s751s/Ojr3u4WY1c3mD/fb5XcmT69VvrQkoWyZ
TD22Sr59nVUJOnF0WWOnTshJWw4KLizxxikUiq9PLn4Yb220L5r7T9WIijS+Cn3Gp8StWSs8eD7P
KaEUrHDrBxX+R17VNriw7xRwoDHzJ5CheN1mibPDEmdipXPhP58qbqKpmtr+6InjCRZ/Ys3Dck1P
bcE9XrIoD8K3XZg92/u6i934PyevBI0kcYdWUiRwASM7cS235KVwdBjHl01t+WBoLcadPHzbBtKy
YGI7s152nMniLAKGP7RMFGDpcjU+diNWX/mLB5JZoIBs7nkHqvG0z/Yl+t6mYxNopcOD/JN28Kdr
RbvUR+FBEx27sk8oWAXvyD3FgdoVjYpB6ho9fLLSA0CiVcvIbEVJLjIECM3FsAEacGnz9T/SAEin
5fT3Pk5u4yx8lhgLWljxsmiFvY86fUQgNvxi/JITlMLw8FwjDVfK6ya/Of0j7izTP6BU7P4dt6hy
woMPEUk1GF8D6vWCu+moWJl/FQ1wWYBqz5ZB6nyTSWoxsPSzYUMsM/hg3+o4xKgKQhfoYetAEaJU
zj1QqWh3MFBH8tlxVEJN0a8FcqlkG5EiqCenfe8y+mrfRk7LMwxzjiEL5iTLDuoS+2cgm8Xl8cZa
BVyMUWhkJPhcdP4lcVWMK0Ci/l4fyDV8rtF06QUqeS3vB3lQyjfhcka666yHGFmV0qO9OWkZyumm
wpcGxQxkpUhuTgTz3d1PWFunv8fYSWv//4tWOE4u2lrKkJvbUMH/xjwm4l/CAavaqQYcvMaPQf3l
A8ETOKVHXEOrNNiORPi3fE3HSjIc6vA6Dggatdq34YETgC4rR0AYnHER8OABaLuZMkPiVYY69nhE
JenY9nllqjFbTqBZ2+LGc6I2E6LX60AV20K2G9vYW7A3xAPKapcVRu5WvVQxqqYy61wI1tl/PDfK
rTKwRrRqUJbKtY6AhSmj6lH+TjwC6ATIJrV+hijhoKXvMJ+5qLfeU0UPzbwh1n8MXVMTCK6lqNnu
LRDcu2iGmw+FS4vmYFEc5afOuirWmtdgZ/2QUiYxeOcpiERmxG7Yi/kztMniInhcWTm+S5I4Aba9
E8Qh3khq90EEKH7AXRYR35oV5VGo6VuqbkRWROIlsK2ejquMzOx51uXHKxckloOBH/meBh5GXvFL
KhJzcLbWSuOVS7VFasnWfHkwWNh7ofzmguKRwav86G7VtiOc/7P3FNyq0Ua0ne4YfeSCCLiw6THq
+H/OEB/6sQUJWYbSgfChHwP9v44/C1SY4yyAPJAysbVHE811MkUJF5EXLzRWR2uoN9x5S1uhlIuj
o/TX2z4XhtswrKtPpjw1OWRZ4pwmmunTSLjimSQBOQNVkP6DGTd8QXUvb3tJDmi9hle4VADPntM9
HRpf7AfQg3h2fxBr04iSTwa0wrlYn4+dW7LKMfhcC3ZsxNwq8jr6q1mF4OXZg7tGz92g0OPHX40+
Mc3wOF7a6TNomwgxSXTRjey9BI9TZS1gkQLZCMi1FQh8H8ZHcaBDFtH7lJzYcv2SLB4vLqw3hl4W
QO6G4W2Lfjn7jZ5fGjOQT4BeK4Pj5Usbk6s8rqkWMHnnvjhDa/CeC673P8e0Ang61XeYYdHmo+4T
vEuiBeOrv/iiMT/mTcaF6orn7NOwX4NmtAYsQk7uejBG/1UbJrSWJsUyBjyoRLFEMEg+NhsYe0ap
tOvOROmKAArNWMAuZxJMuJIQi9WD27EAc2R6Z0ldlpI4QglleyuVdiHafq7G3EcQtKGmvP7zQSjn
YFjBX81yRZ/oJsj9w6AJVvc3JMd66qJ/qWo1RVABp5W0/CObO413iMVCR4CGaxzR5uBBBWgq7dHK
J/A7SupB81ngzYLgZu+gg4O76qUkFYuyaOWRBP/bn17PDAKyw8es8tcYTBSSD/1f8DrnlaR9JZwu
Y0vZOR8ulmxF8sSR6Q+vXFwEEiiKjGpVA+Isl5V6qu9oZwnPCqgpsGXF9n+tqhcokLlZ4/3XywGo
L+SceoDqdAsRE55RdqDLT+Ki4+57ToOsLq2ItALQe88QCdtszAoIhxQhWCQowQp9VmRMc64TP/1X
nJBs6afSnRqHbwHUbVhA7m8YprvToxBkFcU39q/IDnUl8d3eoTZ+c92dEKevML1BK/X1lofC8aie
ficcCI8JrWJV+uiGrD+bxBs48XNebbAK6LHFPkeKB0IgSGWKTVttS0CiHu6RIsY3l8w0G58GGgT7
hNXMzTqLkxuZn3evCZO5x4LRkMW5XIzZsB+MHcEs3NNUHrJMY3qnF2eTn3vZm8sUT4hAbXOi7EbG
xx2yV3y69YGWyy53skwuySNBErqZNJUlmgnDjT2h8LGv/uk4QmBUa4Wk6xClLGqIClzEPuRhiNWM
TDXlkr45y7T83CH+MW6ajUIPuVnUg5gkl/ScERmU8POCcrDsmwni9ta8AQI7DUO67ynn4xdi/15g
5NGDYY7o3xpLThbyqmlWIpvZdafSw74tB1AePH2QOLfQQSsXCzXvUnytbhmLY23iIMfTND4II7tc
kZv+/cTtr/Z8pex7iNc7Wa4OX55SIApJCZEU1EX7wgc8PSh7MlXkWWjqDkaxhFU0QvKPacjBP6pn
SA25fQTjC1MCUwunKSjfRHOl2ZhOk93Tbx20NMn7TJtrJTntUrrafvGL/65NJ8hsQOm7iPM2bitK
zNj10g+lxgQYvKuFw8yCHkBWOt9KLMguJ/sTPHI5d+6NuGcTk4OXUQOHuWMUqMEzDPOMeKdOD8fz
KZrQ9mhaKXyUp+IUqhW0J5UYedEy11FQhCcbzGmPiMRiekeiMQuZlGz20hIAptw57u8CLcZcQq4N
hdmPJscI58gt5C1cr4mHVBaV0NegAlGIYBut6MD5wKpRWEm+nqEgQKoIT3m5bnfDizJ+mtobJTF4
+ZG7FIXjlHbErwWoW3G/XKA8A99qViuBqxNL41RGSJRiWLoHJKghIVzJsgoISfDd3SN4TlgfeXuw
2rHNBXdBYn2eI67osx+EJIVUluQD1WEqwsOJstx0s6S4+pIh3abfDgKA0abNW67rku9h7/VPRbsK
B1L49s5n0nS/FldZL2l5tDUP+OA3zsHW6wEhTTfbzQcvo3BtsrrvkqPzcAQim0BKmVXUSLxLEHMl
OYDqF92nMi4d8QRU7CH3sKS7ZPgYO81PFXZllMXMNB7owxPC8kjH3VYkvXoO/7SWjeurfxO+D22R
/zjr7Ez0vHK709F1LrSkSuo8EazfLkC0rS+p14nalHK88f3nPWXu1o1xbBM62zcUM+knvmT9M2zG
/wFi6ILrbQp1vUuYS/lb3kadH5V1RHRXE3p3riV7NynQnDf00LkXjVwgo2f3MvhymfsI8WhhHXKk
C/DbmqwBpmaVQuIzvvQc921sTfd3mFBScWKkyNdqM/GKvEIoPLpkJIeSIrexwuzgLjm86VEvTYyS
fq5V7tyf2HhoNNmdpqf5M4ThLreiR4jzbPfixHRhdcnsCF/WtjPGPRrlmx9dm+dTVDHZBipGr0Ry
KjhltuydGH74HzTFs+p0uk54HEXwxwBSpY0oSkH8sru7YpMvApen5mPePjBDhzJ8BdQkeiEsbG7M
YDi9Begxdhi1lp8stPyVADGJ/22D3palGRvlyzwds3WsY1dR44trhjveKwYmhUwd7KzXiLzmlisv
yHFffpbRppE3J46GTttQyQMCWgGcZampTXtH28ObhVL8ZiU873EG505Xcpy9ZutJNvMMzxd75K5T
yAY2QPK1oFfwqZEvgUNpNg/GM+andvHDh3wg+viVaHcRTss5ziJOvpvg8i2dLb2gITBm0dL2CodP
s1LfIVxghfFoo0UspSW2VO9EqMa0hd6S1riOZsUqQhRRqgZVOMln/fp+kK+kYPGlWIGqm177FFOm
rECcghWtHEndaM/ylDj+YEZVhsLE4EU8Lvaa9yYo8rGgMMHIFsSk3E65Y+Y+6XmKEtJOB0VW4/rM
PbOc3gt/l5MitLLLwCjH5S5GAu1mXoJ27hc4HFxsIT2b7cRi6r3eNUBMsjs28Yq5u1brh93SqPVq
Lsc6QLYNBAsHVfyv1wZkF1eBSZpp9GzzM3H6bp2VAodV6oUlPzujxR4kEoSGbEXFYbArDPi5NQJw
gqLoI1aTbSkXxcX0GCnByOKzBR08/Tj4LnEjGvgk+bOoXdEw4qCulIcLGgUl9bSVQyGufzVfA9HN
q830kSv/qYf2YOnYqO0opOhbLnwy2YVhypZjnJFMZA77f/hqqWlcdBWO7Or4OSqOBg5VUK2b4Lds
oDcfwYQomXCcwqdyVoTI+5KQ8stDBJ86UelcSQUlZ1Au47QJ2NjaMgx13t2bqdu7o70w1JPpBvtS
Yjx9PPg6APSRVq2zhsW4exgNdyFMu/eCc6FqGivqQgDEnGgSDjicIIXglzYv+PI02X/RWaMW2hZ3
eRSjrqGUb2vHOv6tGhBnJqdP3C1oSOaSeQ3fAEAYvnOfPik2iUdKs6ijTp5dO8Eg0qUDeOudNH13
zLvBT13E45uIELKzc26xvNOVhPBWKrLT71biBYocrltclKBkb+KIWeMKlQQnDocscvlpvDUVhFRI
pcShNq7Si83xRFc7Zfth6uAvUNtV1tPZEaJ+wIVZhY9dsTgjB3jg/HgD9EUqXOfc0bJcKE3/EJqN
qvXL8iNvwHxq5Drr9KH/WvgHFGyWdGiXGsaTJI6YzYiCQK8v/VTz4TcK8v5zemYW5XSWYxBNQOD1
FmQnxXrEJwHRmsfzT9KEqN5RjhvtO25mMQGflO/rdPEgdWAHp0Z6QgfF+AM9Nv2ekcPkmut9w291
ccT20PC09AsFSTUgEfy/nQ4LchnKF4Nco2/AWPhCXF0RQwZt+hlqw3/Jr7TLqjjnV6pnP5D61bIt
Re271rfspPYlpQnUrfHMY2TQvw+ACfQISKcyLLB1T82196qRnJ9pIBAMJb0M9BCnUX0Wvl4FZdcj
L2R2ssE1EMFZODF9LxDT9D9wKO6FatWxvWvB+6Wl56L3jN7aOtcyp8UvKkfdJi5Wrl95hsJQAYiQ
uBJqnnagWfdfvlHR3ItiGx++ZQrxs5FCusgSUCTzGC4zFjbdh/44Nw0ymxbCAGQOAmOTHjhFlYDs
Vnjyv8WppXFhXS3v50dXhbz2bB1IIUKX3UkchN1zGJsMSvu9nBMqpqQxX6Ce2TelZpJTXFzTfjeZ
0WD1Br8D1kHtjeHlcmkVGekCoti3IR+/X0oZYZJ5G8IEoDl42Ekv2ie9ZXV3GFDldnBGnWda8NAn
86cVpcbCpuHAOA+JNfp9GHKT0QnFwfirUpETpa4MbOrsC4llpnuDK6ct4OqOew0IsuPtGNxI+m9t
h0YMmh67v/SY479aC+8Sg+FwRY72GVmSA/2aqMfAee5PAxBcjhIVpUfPgEMs8wkCaP29fnQ5dEf/
EUylsHptBgXjaPqYtcZ0kFF083nXl/Cx/2YQxNBTn71SbaOHpPwZgMgMAGmPt15QDSq1dfrioU8s
ASn8NiUX4dMkA8Y7+avFmBamMzIFqO7eyD6JEU7gZzk/S7YXrZyECY08sDH1Tsyvf5yhpSwzgy34
9AiOL6U8IgEpP6MWLf0XE5ke1hOogdV3pSwBCS/w1AeOjOJ5WWZ7cXMK8N0InkbO4SzDF//L0KEJ
zn4frVSXinMO5Cgfi00IzsxhJr7t/CK+rBmNhA2YwFMVPrY/tQRLvro6luLdf20WmliIp8FXj2Iy
moUGFGOwSPmYbvPdDp6nutduAK29ws3vDvDKz9JRNFUInuo5hVDLRhTWZakARYBijvJyXdi4vBCc
Vj0G137MDMf8uLSalloeEH7z+dxSEr9L9CuAH+WTKwL9mhtTbGIU32x/L+C8NwkubvXsyDnjokSj
XpL+jHIen/0yyAehIBv1fOSyshetES6CLveNG+CGGJ+E0l2cKU9gz7+GBSDLS3ozwKxbmPV82FLv
6RtztFMIfWPQFMMH/ScbijxDnBZKsM9cR97EyG5mke9IACHLhvtbm5imbHIBBfGnC0Bu+hG4sAtn
j0THzLeMFVeMrEWz0RuASfv32UlV6e0Mh3hW82qQEKA7bd0K6lX7PoUUNNyot3sJ9YNnWf2i+0o+
BVwJGG7fuWvmUoYtIFvQPhK06O8ygVyngESVPUVTKOPmU0d5z/+T3o0eXrXQzeNEk4dUUQ+y3PXf
TdkjJvStrGEI2qJgS20mckWx1Ib6NDACZ2lIknfen+6o61lKjpJKQUZP3BGQdaUaL1ifeNv5hP0W
mESp7VgLeinlzbKvJ0qngc2dRnsh+4YdhuAuCnDVjzuRWj5c7EOhtGeF5K6tcZwBH8JxUnCnuVvG
Kuixqc9uZMUGQJLY82ArbXv/sflXvXFWEmZNNqIsW66gcPVfFZxWulLwnCVpqd8Ie1eJuugCha36
fzRQTeWJp+jkjP151wC4oLqL+0VysRmz8HeS7D129Tof3gMRQYQcZY5QzcH4kpTcJwvjoKcmUZle
+XE5kHeKfBwecyiDD1wDvm+OvG/c4xJhhR9zr3TaOBjtR+9vYQV9peMr2EHvsSP92D28l7+eBnsk
pFOkJPZGjRH9Z7jUJvVuCeDeEXcV4eicpAfWQd+ti2JF5hoZm3o7KUAk/VG8lW0hk351vdf3KexT
OQmbvXHDzrfYpNK3os3aRq08rO7uKVLmexSrs6TMGMoNspwmAEq+qoPB3G/3Vv36NJhouTiwY4Zh
FDXU6vV0pYdCJ5jnvG0R1lq8INZOk5yRee0ixfW6y5uYwF50In1f3I7GG1ealtNlpW/Lv8sezN8k
h4ER5lzbgpyOyugMz/IQrOcKu2yxOEyrEucFuyuMXhUH45hg5bDL9QT+aeQpYzqAc2OXYM8U9ldG
xna8HflAQRv8nxO+q3FlcPchBPsXmVebrY3xjuVe9NCf0A1Aa1+ryA2qHxKIcOtTcNVhl9XZmiDk
BocdZSi0W0wicIEqNGAS9oP7t8fHhwHBxcmtNwI+INjuyxYDw5/+X8zXd91gjHF5EMGuhcTy115J
Al9AxCJP2gN+nqSpIvSmji4VrkRfUaFmVfzG9PkQQXKgHpRW8nLucMdjRpvl35YSzdsK2F2aCscQ
HJPVlofgwlrqUYaDSeLyI4KFFyBsg7WlF4r3fzpQSZKRCypeKlg9YMM4tBf9g7FeIwfMo8WTYZTI
8xuRl5Mmp4JC8qP6zDbbNHMRuOr4103ZlGZ76oBzSJnC1ERG3Ntyv/nZAiaHU07OY9FBAXtul62Z
QY/CW/IhC9q7Nh2+AVypC0sXdJIHRyZebnfGubhdugoCv4M6O7gnLDlqcPXMWEQH7/noOP2/NShb
L5GiQDxvEHCzJeHe5jFEcUFy2mGnf2ugsyeKRj62xi8nylpjEIuL8XIK0IsedBVynchUzuIRbS5o
/Sy3Mle9woLl3yu19dGWwvRXJpLmKOL1yKW+vLJW9Ogx+gFm5+Fu5kH7TG+2EB6aujbsnQuMx++e
aVYrNBqHDjzkA71QtR/ICnq6/kFoSS0WB5MwGzrQnQ+C7QxSMwCk6mJcox8KmLGlDmZb5eBfYTcI
DfDBgpODk9GAjyScnTkXlrVcI3YNoQaLLPvNvlv5yISi4XhiTxXLJ04XF7e0+r/wG38+v8vKZsUI
y7wkiRsl1r2LoXoiw/cWSUg/v0GvhHgHAXGVy2oM0Jrcrnq6tbjoeBbuOuBI9yn2BqSvU4nMDed3
CV3QP07AIaAO6a7zSulRPmCrty0sdD3PJD81UuJTcGfspjazISxgAntReazzIZ6Rcd8QYHKbfxjy
ixYALZV+UBtg0hzbdpyUZ8CE6jdIvZSp+E4yaj3bHzjZr7TZB+pQ2PBlJ+oghdq6WuNIKFu7Tq+4
/wRpZIxTDzdUjv004bCSSkGX18diOWKUPFOTMHO7KM1uSn5zfiY2ob+leSLcNPAhMV4Yu4nzWO5/
XwwEJb9NRNNgDY6SY5JADvilehrIv4jYB/bAKFkg+lOZ/sMhkElce+I7jFAHCrygXE+ZPvtkQDLr
PPH9cfYV59E4n2n2BkrngEGTJb4bTQvtbERErlRajQ9+zW5QEiStH+O5spFFKJEkZhKpO7z9AFBC
tDzN5C5yFkc0p2OOdLmelUPFF+7Rvn05U3dqVXiTaYoYl0mZPYL9o98BlWt4D7Rfl6hLHQg8i4eC
Rv1dPLSybGgx6rniePBH5hVwROy6mBmjUWeVzrtsQe2ozDCVF+MXy1awnaRNaWc1hU8fERzoq6+0
BVbfXdpxAzIuR0X1g7TDrQ2iNG3n9PpXxdjzXaVP+sYCtO4HyOrGc5bDXWNIbKGaXEGfdXd/igYD
UZWTxlsuvF3zV4MQRi3JxqEmcgR/gIRcHirMvCMTbFRFbKZtiwRtOAvohBOhuoKZ+OLnc2CLtnLy
qsMoYvH3LDWbcxqi6gGu2cwyGV+kn+Ycqz4pg37CPdi2sBHmuJCx5LMizn/znuXXjmpq+Oe9c3E/
IkPJFUPzg/H9gaA4M1JzGXXthjWWI79ZGeY8GfrsY9LG4H4bBW/GUGP1xI3fZ/g22Kt8IbWEYHBP
QiTwp+dUPII2N/dJMmVC9xICkdZb1xzHheGzhEtckZlG3w2Ll+dO9e+SYYcRSxpqU0dJvJpeOXqS
dHOThjNJcXqAbJr28Zz7uELO1zSj3GszgfVx/qfxStz28gyDIwmGYA0PeFmQTrYHhd4avWwtariI
6w8MmIhSImNq6W965/6ZLz9h4XAaMnO5YhMuk1Y2OX8EamHZZcYjT/2a2IkFVdx9b2h+/d1h1XBp
FHsWkqLwyKsWwfJ1IY3lZxp+y9NLkHrxvyDCSKPjDgW5Gs+xvSR19NZsxSu982AKXWPia/tHEY99
IydK8Atnou7PxW0YJNWUVlx7+69pvUOrOev1m1dj+sRF+AbNFQ8ljwXWdVUEIIEM+CVFbFHo1clY
4vgWGE3Cd9MOXyv5rpIvRsfEagLHZitOVV3FV1WLa7ms4Y8UNUrO1gUEp9WFCIGTN+box69rxc0M
7NOjRnMCDVN4mbRQnZs5mdgLDA0e6wuL3bkmZfVTepDMuiLmTwBvHS+f1GhlCp9Z83RQtapu+CH4
aXu8gD86mI217qUucOq57YX0N7w9ki34crrrobMbewr6j9A+cwNNzVp6vIjDWSfwO76n5MZBjQTs
OR+tCZtQpfoX0595NfxjcijvrJNveX4VDNhkDyZkXj8HuDA/S3xRbly7+4QVZP/714N/kbkPxcas
0bNCvKfcUX4igHS9nyJALwXhehMRWvfdDSUIBt9u9GHHQmWFmHoPd5Bkr4r7G/1xleGfrDggXS/Q
MpSJdCUz3irnorZavlk/BBc88zO4+K8LmdW4RL162eir/MOS8Ee/bGUZWS5uhsR1To82g2T2rwiB
CtnJeaKVX8ETv0M5TjOrCLU/i61fddHil0lEkR0OUhwDeoGR0D1nyE1VPRpWqpZQ/5CKNpPMMYG5
jOxhsLiUuJyKlcGOChJ2IESggROtM/kB06/SBL4i1Zn89P90Nsb/b7A89bQBjw6q5erd75ywYHs8
IqIXCLA4QEsaxZ6EZ8fSVdL3mka1QmY4D3fmiON01L9EuGwgrlsNC69OC2lpn9hONHzFqqgixnTf
VC7689cH7i9fbDk9/4ism/GLX5FpLG3YBK7gOz5JhAWJygdgq+My27rJforxgvM4J37tWMpOZxCC
vPcwTCb0hoy7qKe6fGEuTN29UkGKQmtsiHVN3D34h3r4Y9FLszm+LsB0oPBuKNsvuye2XOkE8hVS
IZ72uAz0gluBwPbSbJjHtbRmUN+6ImfP1JUODGJqb5LRfDpHVk89pqBPkLKapTwRKCdnkBAR5+jg
pyvzAnT7lPerrgM2JWgun5XR1tgsoB5MwmgO5BF9vjvMik+EjceHWTbjHNRmZa/WXvcnvNYJ5qTb
vHBvp2Z3u/GD1ZL3xdyAY2PA6mJlp8d2RKKjVrfTQvFrF/3hwSg60XOsjfxSYVlWUbuDTONYQenK
A+d1wX5+FUpCRBPUXEOhBPFm7d2NMigd+E+5Jf5KYrciQHi8lr+wrI7pjPpKZcA1XQKVv0GCESF4
g5Nys1md7oElsscCqUBGNZZvK6llgMgrOFuIyjhaR123HX70yFawM7i1gShHsaq1OG01L4ZGhGRQ
RkZ/rKLVizMWNSKXdKRf/JnU8Kmu62VU7abn7gnxoZAhkVD1urRfmaPDfHNka7Wd94LXiuevEiPU
faAibSIutVnDuSaU8L0H4jMKbFsQevZ58pDO9JB7hOtpJKxNP0VmCvSBZs8UwzdMFHVXvBMzHn5m
YhqhPNfaUQ9I3fdtvsFkqFcNAun3OmeAnNdJcbDWVqG/vgvYhg0DombKB9ItuDPKI2G1jLqjXLwy
eV3rwPzr91dVytjI4rCXRCFVoT+gg9SIhfZQQxN5UL32HFBqptpOD1IPPKabi/NY/DRdJzUm5WOR
lObliPJNETmw872uAcZOh8odcX9MiOdaPyUrwaNRLUMNAJCypOXZcFv5aB9rBoAuCbUtdmEpFtkE
i9hETFi1OgNFpYhS4htm8u7sJqyQPFQIEerE8XptPo4JSJQM0GOORFAXHhrZkhFe+XLpMz7W5n+0
seEDVl5zPyu00XwUz8nenuWTjVmVHw6RMl72Wi58qjxAEoWeqsPzuW+IU8oNA3zmqLPhtboHsLcQ
C8JACKgdOUZmMj3VT+jsZPL3Ax4l5ZAE4ISXwjj/ZWJLQFViVJ1yRceGFqIaD7mwNJtDL3vdZ+fn
ep1qj65yQjlGGDtEnMjanVPodFg6PurB8N4/C6cpLwCG3KI2inCUxU/fi3a8q9k+sd6+1bx6U6xY
em9fcyw6BKRQmEH0hDMK1kHDL19mqZRdBZXbkziqeTncQcZus8yRjIYOiejG9cx+/oKcrHST4ogK
4UHNzs9sQUgQPIu4bJ3nvxn9kKD7PlPFNYkgwTYhUZnB3fgMlGz9QPCpsEm6vjR+eGBHhuZbMSQC
2T30iPeGb+LCxA9a+KAKl5GDVv3Lk4R1p4d/3ZFY0zHNjUPsflwjfWSYpapCN3xWXF+yJYNIwxr7
FinM+6l6w3xAEnrGyT63oMQ8RSNvhb7kzF8s1VHxCyeuv943JC9hIy0ofHmB1NDzMtCFwVi2Vez0
f1nMXPzYpRMHHvfXoKKxQF1ngfLJ4G7IAvsW8kiQR0IztlGJVr/JqflVFeOO5DsbYjQQCd8E9wmp
WhMuDfo9vpNmyGPhRbYPNchTgxrN/tMuP9Qvvoz9aR2l8av3aIJT8akW99Zne8L2r4TQEAGLEw7U
aFUlXWYWPOjREBLsNbZ7HpTrM8QUdRTGsatxy9iLZ87grgwuhTFeG9Iimb2BS53l8jS43qtZE5UD
4B/6ucOFh8X0Qfbl/DkI8/1z9yaRO2PwHZWHrnsMZH703pductNgOCgHB8iqLEwELptPRhkvwAOO
l5a0T0jNsFgKW86ndnrjhF5U/FQ+lw3QigsW4drNC8DJAI55yFYBAeBhf+FjlTN8Lh6GzxicAeB0
J7q6tYKYG754DU2hRl33n6DChGlRWWIqCN81HmgDx835pwcDtsGzft2WiOGRUfeNfVu4UGdBOWhh
sRPfScIPcIsXu+7k0UHnWb5XImVhB7PR++RgbxuxbiV8gbe1rPAeRXSFKrhewgY8kyZHjASDD66v
lQKAxa8d5cGhN/j7KvSllYXjIMZo9BWE/d/gNtEsuqISKLOykNyf60UF0znhD/Vdpsm9VbZRjQP1
F+l4cVIarOoVrYe6/KoCxHNZZX4Sr7ly8wV5n0vtQwaYtg23ouzSL9Z/tuuG0MRXWxQGLc/TBeUg
MdusdSiaXOK64jQoKnN3sJPX6VKC7Iqg6j6E0hScU0lEUcHpBsyPiOKf6GEDc9Dr0TDBWU00sQFt
YLuhraXpCZw3pDMerP2U7m4J4xJMaQGsKoJc/jBxSB4MLjP3hXguWqTMPHIBKFzGUABgLzcPBYH3
k61Bbj2Yo7SEx82mPgx7BpaMclFho8Tne7YuBVJ1BzG07qJfdUaqgQYg//8KkKbCBdKJ5zL9U9yg
Ud62xTkZX8Hm8u6G8KWlL/3ZLCgxYlKkglp26nKj+7XOZiLDCDyRwq9oWJvJIOTKhtokzQttVAl3
TiAZ4FcfjluERhktX9ZGKDTJbRVUpNMHsRJNjvQo55Rwf6RyFNtm72zlfkJ1py9xZvVIHvVU9akX
sZyzT8TUbFzi1OI5T/Qs0VVS7AiHAI2wihfH6SncIcogSUAhrMs5Bol+V7imgoIB1UZ1rJGU+DlI
FoRWcjgIDOcsKAOjUoKhxwvb2qdUC0+t/FOkfNSkxyAsp2by3HLICLuccm23EmXU7m2BFdeuc6YQ
QlsxBKcd2WkIqj2kBA9e80SH/c9Xpe1dHikYkOcWZyTX4zMHMUvZeIloYl3XKhCpNC/9+oHgWdTY
H2CMJa7xflDtvgkv/e8FTwstg7QjcJSKxTltFBDVX0LoXV52EB0hSTSEM+5U4D3eFM7l1hjhMbsb
swzPaw5C8WT8eQBMDPRw3VfIV/aXIo3M0q8EnPqrRh3qSf9lxdJdIMFi72Il3ftL1edTA8Y9OV7X
OLReBz3pqaq9543FATb3QJXgycF+gizI6tbJZowJt3DSnxStYhnIqCf71Dt8fcNFnuQjF66jjFaS
BP9zKbu6zy1E7jP0WIQ86Lkydx+YzNlrzsx+gCDMzo6LDG64y/1ClrRC1+6ud9m7wj+hRjSZtAPG
K0S9jnpKZ/belhOP3fPLBwvbmeN3NicVO+lNkQyc2BGXnkDhV6Oj6ADQUzWEpCnYArSuiOWowc2w
rekhZT4kSWFMft+wuJVXp+1erS+6qVImLtE167KkfDdGb4O7SGCTe4N3yUhj+IwH77jx8RZ/x5Dv
yr5yCvztihMBTRbtZX290yLGAVAWbY9TS19zxUlmGr3RLR+9eKSBlg+CWQggnxDTsEZz8Xrjzrbz
fu+Tuiv1tf3+bMlLxMnR6z+mFg9A3H9UKn3kgcs/p0NAvdfPLKE96AM7K27YhhEVD6iHeE9CHb21
gHfwRk6eQByc7wqdyV/DbrsPmD2GBxcWBmyhjMfjlVWGQy2CUecLnGCEyyGSSEBOnOTPknDpZ+uR
+lRYIRbq9ULSOemFc+4GkWy6Td5heZOSOPK9Bt89GGpmr1iuj89sXYG9C8eZqJkrH3vvhET1rcws
9Gv98s/+aCg9xOe/rWZN2N32ROZrGOMp7MeHlNYVF1xI7GhZQif6rrW732D0v/WTs83CV3oQ8/7c
09GUzmYvftrLn49r4OTVyekKOzt8+qDgHF4zKTMc1GqlAq1GQAhKKITvvrHzY5dCdYipYT5fJ8Ui
BVlYHRq+d9uXVxTfVqJyeov0W6yRpfH37F0Q8KJr6yNNmW5RxXKCwjVUIfuLZRpUXnFDdwPEfaF4
s/RYmw4mOh0H8fa8NzemwzCvq9nF4fIyvRcQiEKLYfdO78Jtl6MHazJ+mMyYkKbmm9rx+MnqP2UH
LEyzWKj0GcF36x+ELUdQDLtQjSH3ocERPg5igic53XqwhpRsXabtd54AKxLfSYdqIWNsArO/qaP0
PQ03ke/FfuR/+Fa0jrqjKkL7b7jkD2GYOhGn1Ui4NGJIdcbLTZ6U6Of/tqr3a/ZXxmjer4JkOHrw
OlvWA67OEyj/9iM7Z0n+Tb2SOVeKinC/kzN2wKZrdBm/33BNj08iYAj91EzglWKiSLhgiZBpHpVC
H9W4/b1bMg8oD1u+qfkEwABpUaBeUzyDG/GGX44v2RrqWPykwy8JOeLLi7Kd1zgwLs6p44KVq9V3
AQndcUy42KivCm04yFrZMvUcAs2Vl4DkdS0qhRe+G6RTLJ+IIkooXHL0LgUsT/Zsz1mb2LOPYpJm
mjmZGXRx6STJld7NjlyWSZJO3emh/w64Iq1ScodyUAoEf235mOLuwX+sDA4XY/u/8H8IteTmvj2w
pICQukIE09ccDGqvKKZMv9/CFUjjW50BFYAmA+MZxjAvMog9jHUgpZ2Z7MPVIxxJkUXAHvJ4WlBn
OGOWFj1lMGfJ+JQffTiUVMzA8VZ1U5Q0kxc8WcMfn0Gnc6tYYtUyWrMiJVHKQmpwOz3Gmdy1jYIn
AV7FkoH+0vLh+5fU47ys8T+ImSizx9sO1gnthXyPPAGIczxgYcst9sJjS51LXCxXhEErIFIsXhDJ
3OWpF9Ao9zYmBsiIxLvZ3ezdOpuvPH+XFFDnRlbVW+jZPUHpbOp/EPTSfXVbJn6uc3P3f3sw0cNM
q0evR0KBBidFvfieSA2PGzRk+EgV2OgoPG6v4jxLl95tOlcvWbnosgLkv4qaE2DNKHsSpR8gG/Y+
10cieulnMEqowv736DomNTR6e4NYFeVcGLCvmFR7OTnssdJ7VkueCyatE3jWn54OHSXahM+fxYnZ
Ve9xtm30MnuIfo4KGaWh6xD3TwV3jqPZXLFNwf/zECiWJEkG9I/l3n68T1zk+F6u3CpJi2CYYfo3
bVdUO8IK2s4MGrmjGO0QLYv2YOO6DP4rCU9vhk2iizfbg9qwIuOhOgeDWAH6rc2YfvOO8OGPa76M
02wj78PCRp1d0efo4GCfHOLZBO062IM/eHpvk0F8uaM3Gv8WZwF91hoF5lTYcvRpQUyPzr84FQ4v
R8HJMZrFvKCXbGS1hT2drnHt7GPBhW/EHLCjPuP5t3MYEdctvcB9RoAgg+8nUKeQTTGUucvCoQIP
xfy7TfmGkSydPXbZTIwVd/ffyak4XgrbZuFkaVFQ5ObBaHydflifMuQs4ggu0c5XsCYWWXsgZvEn
/V9ifspycZA4W7QD5TArotOKDoht9qNiwOpp11fIQGlZvOE7UTKiMtTftHOPLuppK5xGFeyPKRBh
IyH38VZX0tKic5CLOlAeDzAFVf24JhSOiM0JerkQ6QpUA2N3ZNTmOyWYwY0uhxVOwt9b0vaYMhBh
f6gDuqMq9d49xObQVF1uZOELShkOIdakVcvA7muMnzLS651HjEzkzp31Rl3cdR1iDIE6yYMiJFHR
myTnyh0vc0DnrOVaeeJC8ADS+LY9a+FcSxBGLGtL8+tHkl3PXHcxM/WXPVfUwpwq8g4oVKlyg8oJ
YWQ6hzGVEu99KueHQ45pe3GJrLSG+YakMNHVNc3sG3ycRBjUem46q4VKonapA9CpBnWCmX+LE99P
KupFCvjj4wxu94pvsok6fVOLxxwN46elqJqBYAqW4iusn8H6IozfAs7o7cB1b0BZYBaWIqBYq+13
PwF+QIHWgrpRFwuGpCpTBgSu4liivFbmg6NLSfS8tSbh9wanm79tc7mL0JOXDgKbFCnpfCpJx2n4
E/dhboTJ81xIlYgUis8Hfni1296ZR9c1JvR1Smh30let3QeAcpBU0S/ycskcmBFR2gCV/uB6Irnu
7rTcODp95nJYyeS90FwjT0tLXcnJorV/hX1lC/coXanawX8fQg+1NKvNZUo7f0l8RoN6q/Cc7aiJ
FuagTL1JANm7qaMSA3ILPdFHu2zdvHd3WykTxGpb9qgvi9xgJHiTroSHzMfqXrj+p1E24aKZUt18
QngluCm/jNaUWZU8XxbESjMljUIEMeDrPp5rxoVY1i95fZAeQkocfYWFuDl2Wd8Fb3gQ6XP4+Shn
vB42RZRlZlZYsDVw7SGcy1yQNTxvZieJ0Nn4E+9IScGX/OZWFePVFjeDgHeRgI+bb87xUQp/Zbhi
2jCibcmyHHU39jZ8rwa6j3rVRpfTbo/IHlsj1laLk+jfjxUkyGlU9Es7n/ANp1l45zqxvMmyXDF1
z2IdxP0ToxsWiDNMfj28hamCNyD4Ze+WXvuUpbAzWmnQR9iZHjEtqTkehin4VbEe4YZhiHvKyCCk
XOxQci8YHjZG7HnYHDgjjKHN8p2fIV1rHlWq+wqx6JqyCJkxpt97PZkOv8RaYcQ38EdKBur1rMI5
bxZz6LB0yyBSXDg9/YJkLCI5oCB2REsDRYybHp0MNxQx+TEUj9C73i8QwPWblX/Cm0YHCEGGL/5Q
0AbwxQm/5phMpiXF5mXC/Q3cMq9CrmQ+LtqWRIX6my0w/Yb/EgwjITbFBTLidxI9ZLtp5vq1S2gS
hK7puvu7W0vCEhEqb+vfz0lqntl4I2K/U9SFprAx+xksshRgGTcZC5qycJBuBbMWIN5bfa1l4jT1
XGHDkM0RSfU4pjut5fDDUbNsNenNTlB5jvFCKX/Av0wwJVFa1O8iEI6I6knNfhN5iSZBo+eliU2f
UsH3mPhDYlQoFbcvpjt5uMDxy1Tw8IHb5MZ8gcaVaGCsmsgHi9gaDTwfKtXxSnPpV5MKKdil8v30
1cawjP5KFRIatscue3FTk3O7bFQIb+GbbSGrBCoSz2hWJ+3DNDosTO4PBr9kfif4hsL91h52K6gN
DsHCohnTz0108IkAxXe7+2Eu3ZwRL9TCslP2BF4X+Osinxj174SHGwCwh5x4VOQtFuUL20W7Efn2
2Z8RU/MhvxjNUYOyBNY8wVvQ+qbZR3CYahLWg4JDE8+xegBi9tACEoW5dpErRIcpKOWpcDLoTuMf
9cT0ihsC63El2CFGVQg99PyLZpBDFpCvr7yUjAZihbJevIA61oMLyinJu8EzP3WRCgFFy37aoD0f
fL+6rTKZeX1a5/IlUmxjROWBa4HhiJDxVdsf4IOIDh9spZ0ZBYyBtewfEXr1aq16gkT81rYu5vB1
U9q+sUxazCrTBFiplZI0o7diBqtPUgLpkiFaf8hZUPPkDyfv1F+JJJUYkeM28aJ6MYyC2DvPeP6a
Si//WIrOvNE4oleA8zdO5+Lb0Ke8a6QuOCTeAVu2KiGmrugjqeERDaIVjDKJeXK/5K4OWQdL3BO3
UOVP8jxihWY4B8f1TwBUO/V1j/UKlssHSN6vQaMl1yOczZllGo45zZt3OW/HySwXTMgGcdy1nXZO
/+94t9e+nub6U9I60UGWf9rqlB0XB9YLbEpTodt9bVbPt/w/u4LHshkdsNjN2ieCbr4K53g4QoFd
0kkgUeO6HYMS78qRuPU8fyXZSCAts+pQla1toWdgd2OeR03BHVOJLQkbQH1AUu+pFbKZ5UWQS985
vMuPswoZ16g/04TnQb9TrlEw2KFjrBWR4RnKUo+JV/CFRbGxpi1etYe3k+goCsxf/Ft+shWOS3ye
25LMt1lmB6Ntr4bHiq9whwyobrUe44Jd1bQKdgUXh4bTtd32F7hH4uXgwONEy9zvhwFbXgNyO5U2
RURZ5Vu3EsWcd7Qi38eszQ7DTogUz0+s9yjd4heM7D9v4CNzzbBRHZW3ZqEokXwAMXV0Q1RfsZ0X
04Bs7GLv9ZEfl+G7QiM27GP5XXlTTt6xAKbFPi+VFKZt8Ro48d5I+1yt1TZXCp3ni/vdHvxztMGC
+2elxGENwa4aCcCeBoAbaiTJMroeE0gw6jt7kQ+HEa8Rv+k5zgFxwFyld6lBzm6sx0JzC/kG5yAy
yffeNQO02DAp/euFyycWzi4GWP5Pkaa8RQQy9UJgXmc0+Fao4raRoyxYyzbSzVvX4dJlufW9QFGR
s1Ee3yMG06P6iXPQ0ur80m6Bgyf3g9Em+9r9wkWEw7bityvb7EECMIx2Lq8kp25IblxN5/CiwLpz
jVLHYHbfCcRHr6aTjLv5W2e9pDr+9Ly9S2/ljsvGzjq3z150yQt1KtWqAvfMs21UrjwBSYptGmvf
JV5zJ+iohXmau3dxoAt+diNfIOy3aF6CkzKmqxBn75JzzM7BrueqDk2HMBUY+KG2vthTHlmuDJZI
8TIGPFQ27LFWBFy8f60WKh//rg5VPYSNe/VxT54i9efds126kjArlfCU/Vg3uaGQtuAyNByynbWG
26Zscm7YXtS5rcShycn//5l6Bi2Cy5raTHFUpqjkh2oiIwl2KO4qrkKqwuh+nlpAq65zUNLp3aBJ
ncjxOdttRmnAhFem5Xb6ESv/29eqplpwTqqj8TPINstLFKN1EbEoS8QWLuy6vps8h3LCkxsflkv5
BNI6sDJG6hVfeg1AXaZiETNycBcFwJKPN9V4ZDYmOK6q7AU8PerOGE9m2qdWE74u2tW8qdm7zWyg
j0xUKR1uLcs6qyvIsMW/JkAHHL6h29sMyLbVdVsQvXtAc6BVFveZzXECkg9FdbMuBWbMSNLflJTv
n4Wpk5M1v0la+EHH5y4BaCVl5plcWfAl6JIWe+4l2ew6VYQcsBNOJh9qU+4jYuc0wGFh2i7X3OWd
Q78pl3gAvnDNg3EOie8eSbp1Fi7h2TGissgny5N1pVUpLwPu2V+yzezidRLo2Fw+4FcsteCxitoW
Ylmw5+ZPm0KFB4XRxHR6ysHR5XJs2JIxem30aRHZzuGuPzZhxYtpZK7JYv2H6f7BOwBKXxJ33l+v
WzJMoAsVYOSUROUw3KLlM16jTIac4COmyc7gaCNxvMCFVnpRPYRoDq+XnAr2aras7scdq7NFL682
BAUnr7dCXUYHuz1I7TiVSvGbFBlXLqAZHD9tmFhgF5lbLUxlv+QVfEi/Od54BBOuGDlXb0XJQp/0
16DTqjS+dQbiYr+YcVz0/qo/pK/ngi2XbPlNrDnIlT3/LDXUNP+i9R52Q84/GAZS+F7IWQKAiQUY
K5EJPl4YBBOc6NcuZzEKsMdTzjHuVEFzafB2Z+paUvVP7oEWYli+ODDlKxI/DzU6rbFs00aFKTM5
RnIkXewLm/EHPHvDtcahAyhD6BAQbjnff88+HtAFqrrqqpWEo8TqnvM0lusxS87e5IgYdQAbLGpv
WE7n1eLjsABTmchslNmtlf8KFxCs6lojIFRxxzU0LZWSI4zwrpW+wgU4OXuVw0sgNcKXEPg/ADi6
sPX6JOsfWXTfBit5coR2gzhzYNl4M2OG84Ze8WZat8gGSFRVXOzJKnMePACQmh/tSjZ6/YPg4R9p
gFsdcs9ggYqGcyLJr46m3WLJHFuWaDkUUtwzlSDvAlSBdv2pFuaBtVd2eBHrQfXYPGur5RSGupJG
AfWpHXTX6vCC6uiJ++Q/wdUjxEhmup7ErjiKsWp1bzODj/dvPqp5pCeVCUA3QnI3lesRp/+M9ykY
ZZL1Q1C71pP9ZI3xlJZYo8+6UG3QGhRcazZ0AHAg83AQpZrjR0XQikRmaqDyGXB0AJtplNn+qePY
qRbQ561ts9Du+AWfpxPFOPAke59SlF3deeYmq77uaAZqHS1JJ0USLj2kBpN32zbxsG9Je8WyiBKN
2Qe9Ogb+LMbD5hkQIVQC1S0y9+mQ6VupCRrDZgCudtN5oPKAjp7AgPAKZROlFvuz6fRSgN/9zQ1R
uFHs4Njfrn19+jhZUXNxalqhdoboA7ALRI/D+rqiiCVMgNhWBL9zJvs00OQ8OeCuZVgVwaI9yDcX
FDJAw7blR7KCFP6pK0Ub5nF7JxWhmJ+ADi/jH51aQsaPDyyeFSN60yBXCq2VKfDdC0U6p/32uSTu
o2ZFuI7XqaK5eSBDnZmdpU2wjMuYNZDsFuOCCqkV3OY6qs9VIOlOCU2thXfesoLlXIFjSyeFvjv5
GtcFxV6F5x5Don246v3Fb6mP5v52BCNkHUZpbrpm1PoHBtUV7NYwEIym2VQPOdx6lwYCivPIzulT
6WAJLEOP/LVwM2Ko2zR/64Dvc4sOw4cOq2Dxfq5A+jY+5GABsPEZxrkixGIEWuUHF30KJBT9qxNq
k9vAgyAW1Sz2WxME7MJctCLS/+t64MR8MPZG3128+T4MOXqqRzulD+23nQUMLi+nUrgy9JVBctfI
9aQvVN0/Lb7PsO7cS63upprJKATNSOGJnKhpdS/ORz4AtF2th4dbI1fQMksGxrvHTP7hUbdQIByM
LsNspLY21iErJJpwV6jQ5BZaPoDLRSvnnyCpLG7pBxypujoC2qf3Q9aJ39u4uEoYkB53rspArrxw
+wPJUXw7v8XvknWJfpFifwcEJs89kCUQpXYtrRDc+GWztxXOmIcq8GCYyotvqqgqJGFH2Ayf854h
7y+q9DyZ8bqM0DZyI2oD65gr0SHpMTREawAGj2RLFoMQixiZnO90NaoDz6VtggGFuvM+OBUj/wgA
msDIJ4gPXYMr+Nh6C4t3ORoxmGKFTZWy5YRRCOX8CMQMgLoTzp49SQvMRCsq4Sn41CfNoK+qzHtW
39DEoniNQ1ObitMFWXfLeULpDHCpHhIOHBA8Ay/cfZSH28rzoeLHfiTbdAN3OjcB/EtuOBhDWbQl
Vn96BG8e0lzcLmy0EurAZIY8fkts5+DHNvE5ovua2GcqJcwzxady0jk74EAdE863/JQRLZ1jD0rI
6sxkRM/v2+uo48sVF0DqkCLG3U4xLHJ092Omce+BTrYr9RwnGa9i4RCftzf66PHRxWZntfKvfgK+
SHZ2yWSp2yJEzDy8cuJAq0C1ZaFmQKxF43QNRvjl+rMvG+NXLI1LrUgMMp6JnSkIlGP6q2+KLs2N
U/FUecxWEr1PRbxNGO2gJUaNtT/ZHsoYjvv+JHWIXhhN674rhbz9/04PZNNJIyitLzO09ABWBO1F
Bbd08jskdDDoylHNY8AG9FfVi9k+iTrNyMLzigxEO8HCTuwsF2wWTCkq9S46J4d5kAhNfnGFmyuU
8KfORl/LX05g1fF0zATZRxKQkCTIrFgp67D81LSxyXQlrrK/20/JbpjSPdRMFh2lDLAc/WZCd9Ri
maTh5+hZWAVSBCdxpWl6bD+soJpKtdILKeaKF14sM8Qq9KJL9ZhYSe8C4KUK6jywpzshgc5YOYDT
3SwDMZk2xSrzQGFbcgYePsleXCeDVq8kFf/mMjR/B2YJ6hTKhzC5IPJdxJdQCzpEqdjZYO8XmQt6
ffc6kzCJoZkqlpKkasLm2/PLY2Ha5CrbbE4IfyJMgBQO2mwVWW1b74NjFtOgOBbR2nXcX/HphCDJ
D0yRszxiCHvuuImSQXfHRWyWx9vqLU2+JWraQVk10eBbdvasEKoBmqFL1dTZQXOJ/Dnmb+37e/ur
KktlqyNfIvWNuGL8fv+Kbn30T4WZK1Zt6DDlqmLNuHWJCQpdcfsUeZlogEY7tO2+yTwRuM2QuJsI
qGlUD4rMa+rNToByvp+kQEzR713jdlmjbqQJjp0tn1KWhJXGX4BQIIkFtMzcRRJPi26J5/dFCsxZ
A1n8T5BZUfrtlTq87m4b4u+M63d0DH8AehbiQoODvjHR0AMUZ5MHSptUdsKIp1x7E6jJnW9Iyrah
2WMVsx/AEQb3NTBnka/EIKFXouHuM+TjArdOzaGOnGTN00s2xU4vQyQtl6ro+hP34NtiTRs2FKSA
71UPH5Itkw/d/NURrmBciV+XDU9RCfSrD1IixZOVJHtZEqZrpzqACc0ddbXUYFoUXxFiKsO6D2Ew
Pbrp1iDf2BymhueYO63CR6wYHKPswnTB3l8DRhYtzV27PyDDHrTJTzryZzizoUB2Z+93i7Hz69X7
fWi5PsABgxV7UESjGVonslcg2niDxFwJilBmrKrH01bcKs86QLIx+2OaXIowt/Zax6KUTKCNKlPL
SaeOp5/wH7ZIOOjxnbGNsaOSyc9Mmq/dKETljj2B67ym5yZyCWhGPb1PCfL/bZUYmemBAGRlL64C
I7i4nhuLGkdAcxrf8lLWh+nQjR514Hl9XfUNh125zV6yiCSVCJuUqKgUHW4bAhwPr7S4kOmUTTSO
uvHElsufZ+YkpOwqVipMkYdEycrrsvbqadvcg/y7vSpIRIkLneuvwqGuzfwC8pLqBoDUzz5QrV66
rKmgRTWZ+nQ+6LHr5IF8/xir3KLZZhQ7G3jOTqAlpLWVJcQx7FKRpziPcJUDnyYx0E2yMf6JIbxk
vdM9zOwW0IWS6e2J3mWiidQSiDIqRD9goEY7YDalx4g+IaKPMvno6vfrWxatP9O7clT0UGizUZ94
MaTQpcynMcqd4pkWsUqQvxajqPtJvBF8jEb2dgavzTj/veAA8Di9zJhxWb/m4vgKIKC9IMOIQW5i
NXEFnnH69AgkaHl3uMbz+xHvqjHYPSibSBpi2yZlWBs/W0ea+3g+8HkmqHRDbnPiVWDCVqMMUQTG
CuQiZKkSfRkpZ+wss0dZBikvsK8BIDw1le7L/OWjA7NLHI4ALsoQdsQ7FODbDXO9wjHGcsRRLJFo
UB4U7w0OAwKpYJBUIgZBAGP+44vRD8aupAGvk1BQWf3PEpVLYb5KuJmp7XKNo8R5mklawmx4fOXB
WJbY92RpVFaQ+QCSOYohb/5m4i/mxiYMTek1F9t+vaNUdo3rQg8GSrueMGaLjLEE7rmzVlgMo/K6
heJxu3u5EMQiqYnpovaecMFApE6ZGeeDWds3RbdZGr4EL6zkBkw4Io9BwcU2DdFiA/1BL76aqX9h
o/f3OTN9EZ3p6KaixJg/QcuZ2u5waBsxjPxSo/Izqt6JVn8JKqe4lKkzO5sck4NhQGmma59sDEJk
xqd2M5+AWYjsJmzo7lwmv5tbe9NyGIqhkRbx9K7ZPMgy/F22D8dOf3HYOH/pu/RDgK36kX6qkDfI
KbJyUyjZ08TKbEIsPnlLhv0lGLfZoCVK29S5rVM2Xx10HIZbJh5Zo3Wulk+mhIJAHA5LSn3wUfhg
OzS+sg2S6zSTSfUX0A/3tLzWEZww36XfuXEYXyQdfl0jgmqF15q654FM12lr1ZP/IlEwJyWMA9Oo
UOgqU/9QkSrDPfQraQ54WCAq7AFz7nIrIM5A6+OH9tnZADKoyTJPWmJJY2+ZKDJNMuSRq7yNh+1M
qPFb9N1FAmDCboWxsm+1HQbeQBT8bOLkRn8Om3C2P1A2n7UmPvPRX6FH8lBoZPlZ3R3upU5KzEwh
W2w4VG4Pl/UEzsXnhqSl180nTbzFJ1c1I3SddudJvNiMQZOVe+onYUu+slL0MfuBLf0ze6weX6yw
FMD8eCKQBdiIDjDxJL8ckbela2SXLVmYMq/20X2nw56UXlRRUkh2gY99m8urQl+yZSLfnEgFbEkn
nYlxXpWycwkfQytb1g6xTQ6MZCujG8u3t2UtUaYrXZo3NgnNdN49xRnmK6t+8gbOg8QMmzaUMy1h
6m+hT1NNnyscAt8ZezcAbV4XJeQSkg6KrFGnhNCJD0smgaeOWim+1QPhLTDel1ApXVRyDBB4TF8m
ABJL+x5rgv9S5jOHYh4yipmv2ZolyUzJP9tA72H/5mM8j1zrFC4Cg+1ycvjHCy6AxBJ95ULMSzLc
qRPh78EZ+/WVZJW/mkGe+r7JxciTNvJNadffmbEFQqjmQ3n08H+8dN6o0Xq5efjZYQF6p0BZiPSH
4ajcN809juQKy9Pr85Dy8g1HrCJ1LZRiBfCrSEtLbNe5GG8CKAEjOuZ/uEFO2layiN+LP5TgwNbn
y4PI9eWs2Y8O1XHyPy5P6kLodqlGNMe96oqJ0rWco6WSECmhjyedg2qL0kDav83u621SZIUPfIMi
oEb3el2WsMb3duagIuFkALUHoBTSktgd2icTtjWyd1YyhQct0ocbog2fkE2ATA3ynIjycb7KpbG5
0tP+U5/PqR1iokvUwbQN27SbsSaS8zc9lsqFo+815d29WsOvowiLNLj1miKp717Cmzdr6+/vO67t
k8jpxbV0EF1zQ8vyOEd5GSbSMq7c5fgeK9lpiQs4T16nk5mudAd1S3Je821lHk/wmnVL56xznn9J
8ccIh6Nz8tN4Mva1R03UexZxNrrfUNy5pbxqEo5/4dDhxrBOEBa8vhlmILOU5B/LUiGKO2pZjXWg
7dv2PUapz+dTEQB4NqYD+KBsm9kpNgil8F1C8AyH9+s1b+StpHB7ZtR7Z0jDeLtPiRa8IeBpqPSb
VN+WZxZYKAI9WU9iRAWe9cRM4spH3+AhbzJq71HA6DoC0JyYDQ7c5xHEa/f3GRiQviPygzF1kYkF
BsZUvSUhL4I6dqr91bBbXMOolUOXJD4flv1FBx4xU71YTD4y7WDhY4xkMRV+25sFDl4ryqL689W1
YDToH1zHt1cBDIZ6c0BTF4WMYL0Ey2X92YJQil02G7nC+EnuXzJROKBIlqvEE2+7xNIeKVsgGPcg
+EuYBEHkIF2m1NTg150beSOBaUV/bBZDIws2l080auO6JBCQD+4zWRg7UWSE2TyQrKq3vqODA71n
+okNY3lFnf+73I1BQP5r08nVhb7nI4xIyDNpFvTTKxt378Jegc1USBaSEEj4H9OPMsB1BDp1gn8Y
A+IUmPNMm2BjzyGT6hD5sQkOfHCnm3H4NH3Ryl9HU9qHzVILJwLzbO0Zz+2qxx7yMG8aNIgcp/hm
5Ii1nVq8vEXW4tQzwScnzUlT6v1AF5WaaXyT6vNHAvUgOOoGzer6N2WclRou4MV+FLLRnXduYHEc
EDIOvsMSG4l9V9veHmB+L75bEUZGE84b2OyB6iEuzaWtU1Tsytn4VspadK0gj47jT6WA7JZcJO+2
PHuYVvDhxuD92a2OGhDYpOG4RnWddT0CbYkUi/P6aA7cgojfrxSt4VhjgV1xO79tYpHXzumQufRB
TdWZqxp69bPnipdNO4qYj81KYqJnN54J2TTAUQF5Dt6oNMGVRXMf6Bj3FJUwrUXWQwte/2tG4Q/+
EnMp4qvyhL5qAG1/shWSJAY9OATplLIDwKezzt5YQkd66V+45M8cQS0d9mV2kBX9HOkz0gF31k8L
zQh9CW6KyITcW7RY1RjmIksrO36Jl0kTMnUdaEDpC0rUht7KYUWYLhHZj3puxxziIXnKY23MIqzR
ot7uVQR3I8grxNX1Ny7BFQaqp/EESt08S5jetidhH7hUOkukU0pcOdjjKUgXYb10Arlif6HfL0w6
MJEe1zyGYUq1oi/xObetd7Eue9vul6XmelLNxvEI2Ub9SLeafozXxndxmN6NtYdAMgIii8oLxmsI
KKOn1sq5T6I08w7B1YGZ2jMbap6hoxubleiaCcrq6dJTEsqLV1dD3gciNr/8esV9t7XIqyCyPNQ1
XSY8Cf8qZJkPd22I4lkr6q3KGcNEH/VLg8FQRZclhUzAqvq/89tmWfC60xxfcS3Y28q92dSG1VEk
9dT/Kce6QQGAKtdk8ZqfsmkUc0llMMWByLaLwZYWc0aRVxxApDDko+hG87fi+h09iStiBGwevmto
ABCaTQtc0ce8xG4CCqEJlNCgfrzdOMO7RwgUiYhlrXnVdvFUyVXjFAaFHzWn7+eE3Mo2WZ7/tI08
L7qFiAD4uM8EDVTWoiwsL7/T7uDjixxaR99IZjVmUmT/eBwXki0AuRgKNCWhHdbBXRyOLN8ViYRQ
/O/hztglCIDOAbJ9LW+zZYHu2ceoGAnlNqNrVexhwWuh6z7gopTFXGKoENXgbYipCDFxt+CLxSdb
DeBO/WoVhu5QXJ3t4ShWaV+jW3jEHCXaLmdlYNmNh7roMTzzLJD1K9KWyJvcqCGE9Fl/VcwDENd3
je0KOVbCVTv+95d/cHUTTqICMW077lCW1VQhdNIYLyvGeDsYUu8Q7hLdp8BCAsi563QTGSNRT5hT
xCljt41SZJ8Ro+pxVeiD2o0ViIydLQxTk0Mxkb3Ke7p3OrVLOKXcXkGe+Gb/pXG7BmX3jVWTgYkE
x107i1Fk/pATku/xBUFOLNhH7p/Kf25bJ6FhXMUW/7gJDkPcXOHe/lgajm1RBdZSwbpeYzkgXw3N
b8AsMqjoLmIEGt+pWJ+KSHBQPAFnbHL16maDQ4LceAlGEMM7bFL6YTNDJyY1PO1aoCv1cQj+u1jW
nhL1fEYWYrDUUlx3ML0Nc0Jx1BisY1FMrKJApxm6UTmrO1t3jaO43GrfoDzPaZs/Po67MOiKYo72
h3aCCMMuae9w+0RUUr2VAcQvI0bMJOPXakHEiUycz9xWOG9zZ0OyeFngZuI57BuwSQ/E1aSLrJbJ
bZakAouhGqe92VISaCIrMRVlR8CWI33QgwrsWt9GUDzZJg/dgYPcRUuOMGEaRrz2ZFQp/ltFH/Tw
tU2lyTIrTNYYIaDUnGu679FO5zKXUqTeXotwvTYzvQrnadfpI77qJWG5t/BpII/sIab7usibQIyw
ZXnhOA/6SS+GxC2ZLrJdKUMYGX3RxixhWEt5voamGdZVX4rE47iT9CBkaVCsiF/V5KBbHclTJYrC
G07SZj+vzdOMT3ZoaBAPn3pLiYsN6RIOe114Ht06c20Yx1cfsdQpIm0lF6UXCK49v6JiOkl+3wfo
ayr/FH928ZhnwE7e3qOdIfWOcwEMGeU0fqLeYZnCElLJB7TOgtPjn3TrkPnKS2Pvq/QDyhB/Z8xH
nsnz0Ott0YBh+EQ/4jm1vgS7geL7c0slRQJnfXrhPIN/SCbApZTlQJqbIBx4PcCl1Win1bGk1m1o
Y2ZxbrvCZBIB+051vKDYM8wWPRjnL2QMbgIbT7oflPdeQmNkZX0HluG8qmDjBa5kIm8qwVES09E8
n6jCdrc6VK6GwLTtHBmeApm9qF/Du65DbJOIh4B9pcDwFK0u3n1HaDsP5Dna0NV6oaScGNDd3ccW
2wL7E9eCHS/B4S5bqQ7Pur/63kVffzRczV3Dov+rVppDVhaITyWIa+08Gua0lHNqj9iipVBkwWC8
RKLTekKTkoDnKpR8Y2MQjIbnkKdqm96+8Y3ujqlx4unzXtClqdEnfsEuGy/W9D8Y5VOcATRdRfS7
ElnxpJK9DDaoj1RlAEmx0TE5+RcxphHOKyUQOvDPKBKddJ6VtVCiv8U91J3MXLvCKXaEQsSsC69/
4ObsIg4FhtCpR7FDBEn0PScrG+eBG9wGT5JuhlDjsKF2JctQFQK0O/J9YoYk8e/CnTdKH8BNc4l6
1Pv2k3Hu/pxo2V9CMKu8nsNnv28L4YbJ8qj38SZWwXRe0i1TR9OHHGcVH4A829Cj7p8eAOluSzGt
f3He6Q8bxfQL3MApYwVJXHuxkWopLGMl8HNr4LZAbyew8LLJdmxbhAUrda5fgwfERjMGqXm0T2ds
65vv/suxckKSxPR+Jtj42zwmw37OCMcJUcPML6nFwXRu+ZSegk7/nXqxTyesoqVMwoRZdqV9fjk4
oKe3XUeEQoJRSr8qaoVySYeP7Q9ngsqBhcYzRsJIjov+nSescCJjGnEzwAMlMTEF6CJZY0IDvZdk
3A3G45v7Pmj9VNce3bHZyjtQsbI6abNog7URVeDmTeEGQ8KpErDlUHoj+ySCaATLMocSN/F1irP2
oej1/vrP09iS3Zqk+31RXqQLuh3yg2/BbEGDsUIJkWOjfJqCBG88vSf5HnicTvCJYhOC6dYSvxxk
eXat8eS5u3m+OynnJnMctvWjbxbtt5U+b4j7FQFd91R9f3PEnof/3QPDdBFtsphzBvDBDYaTgVzp
aR2vdwB4KY8/sc/R21mpj+oJvKce6Nnb1wqqav+1995lu4STTeHyb2neS04WXxUQo37tDhW9eR5J
XS2HQu58g2ExZx56VPttwq4JayRkyu8nFru0Fhki6z0y1KiEXJhSOPVeyAiXE1NjqOY7iXURa+wn
vZBlSamLLblvLg4s72AyedBO3/g6MIuhXZDSzicYDlvuzfn+5m/1ay4zXP6Mb/LIVrOTyVtcWMFc
PkMcPz4mZIGFguFczcrH93MKx949RTaU8bvcBKOzLBR4mzQZt7wosHK2PGMRIk1473RQyNXbV0i8
tMUQ1SPiicic8Fy97jOjDi4DAo3nNqnAdub0nr3QYYwjUOCwAU98pGF3MIEeUYK4phfJq5Mijywt
V6zI8OAP9qfhoXVdAxgxe4E+pahmJn7hzzdzfb8zIdhRcBZ51a6B0DDsO379rmSJvK/6lh+pVmpT
XMhHuopq8cABJzXJ2KrXsE5Xh/rmscuxSAGXNQZKe1l8ZJnxJ1V1SvWjVgCNMiTRDKREpQTMvzls
Xz01CCoO66V7SK02+pNDEpLk2Q4BZG2OKzTdNwNGHqnOxDrIbdkIVJm3mS7NTy+1j5Rs7THSSgii
aB/QhMkuwCPEUmuoSwKcT7kyWZlMzGKdCj4jXAgfpTog8R5NLFA3j6PSlvr1MBw8MWQ2cC/D9JXB
heq9yWpetbJsRy+gd0OG4phvEGoH/1BCBmXZ2vyeWCcb1lsiN11B+B+ze02Vbd+xvZp1SuecOTtZ
0XYxmEuQgdQNieW2/vzpWr9z5yRGyn3FClxe6h4w/Jktpx76YlhzSXbPdJgx7V9L3PJ1Mg48kDyG
c+eFm+YoFlPAPPHZ4HbtMxmRmq0I7mKXc8whTBgNB3zD/FE7k0qBmSdYhtdC3kJ/apcxdN/X6K9y
XewkdhcFPMHP68XBBx86lY58N5CPXKhGoz7nCuOeVpGCgtr8rjHGwpfiJudtryYhf0bzZhTJHcdg
TMMEUwa9DYF36hRCs8eUPCcoJ+WUh9Lv7gc2XzMiJfahVzGjCjG20M38Kzj509X2M1mYYCzgCEDg
gvhm5M6lHI8UaegQTeeQcSGAKDe31i/X6SRI1R7fQY2b3yfCoUv49hYzIdWUSKFP6wdNduFb0CBf
hEaHtOElKwyEuDvz0Nw3ZjUmvEab7umREp8KTHn+uGMKPi8xShmukiEJM2AwIsfOZlZRb5QiV/8N
f2qv8psv4xnnCs1qKUOB43Zcor4ZGguSdBHZ6YQva6OhChxKNNQsTqo9nI0RaiEW+7WrAWaRBx9N
g49VYGreaY6pXp+ZaKYKfpe2333gX6IvxfpR6U595gHLp4eeThbSQnyKE/KuV99goc1JW58G1AWW
8Ie6Ep7U1bR60KBiJ108uhqjH0gYW2x1WEl70qYo/oHJSHbvY0F32bTOH5PJLXdbCxmArbxYClvn
NOQTxBcacpUYrV0Zpd4mH7XxOJlB0BYAsT9YA2uNCMxPNwutjPxNQcfvMSVSRZJrRgk4t3NYKjJx
tPslSBMASrj4GIH6b0JyYnVRTFkSSiK0NfuJdxKbWPny//nv3ICfS+K2r8LBsKDMQe8RXQIrnejL
8zYvpsyP6A+764dCNfSFXh/IXnlmTKyGX0K7V7UFly3TwfkOOubHDRu+vOOtLp42Nf8VS2pIxljL
QRsV/vqsv1A6QvCKBT6V3rjIYjCuRH1XxkTSY3OF33QYxEH19hLamDu6PEpwRSuZcn4f4bHY428z
0nn7/XiPrckdyRPsx9raDCjLkov3O+1bfmoJqggfwTKDE4N9O351/V0xvfSmjo7FFW9FNyeauuRY
fmiOXJYAJkbJresAfIcW/N6wDM0VBFMC3KZzEQZvM0SA/b0El4+cm1hAyx5Gyfylh4R3VcW5e+wz
ibkfuGCo/pc8zgzoSD/efq7ODdBdWy6P9nVAxKQshO7GS+sQ2KnMeJwqRzQ15Qx6m8KCqktxsemG
TQ0EbBk+G5xaXYRM71uIthNHleqAc6j5ACmjppaHb/ySRvkPUOInB5TM/GsGjO2rSk3bA1juKref
XiOvbaSWk+K2SoKmWzlZxnYdTYDB7xG6TEmDg8g2vykk1PVI/FntBdgTI9NW0dfi9Ip8/bEdcaoR
p3A86krhSK4cslcfxihj7iNXFmXDCZMHu1aDZ2K2wOmyPIhfIhp1bwhjaizyLFL07S8fh0dk/lQn
p5+UCNAuFIIomyMoFJHAXbq9tslgWm99P5hKBDgeBZeXYqc1p8g4kvvtsLz0SFuFwqEMYlsiz5wE
XYUbpwKzN4byzjtlrXRvMeCi+CrTcyeAt1w3pgoUvw2ABxVGHHm8FLHC8YTmfhIwXiSUeU7AxdYv
4rEJ0clt3OCPnnGilofdxGiykD9OdzTBsrJLUu3f0wCK+XZ9mijsDWhNDxj2pKmBuRGtXyhjEVfN
FnNw/l0zy01yUVvLRQ34LVH5SG4giEWrSg9bkE5MQlMl+cg+cyZygG0IRJIznuVoHna4v0WfD9AB
o9yDV68TYO9jhfKa02egvhYmTvlsFjblwVcghdO1JxKInuXxs3JglVA1r0ClqaGTb+Ye2oLttU2k
fEsFL7qZI2DCJtiB3o9XL1Q/X/7ydk5t8e9NNHKdpi1RCAAu6EqNXlshRn8XRaM3QeWvvdwHNTLF
TQjPlzHx1VGIm/qrlHFXuIKJlnGvhkqFKjFdOAmLTybZDnqgghRMjyaqxNnh9S2dllirRxnWJUfA
76nD8S/Mm9dZARfzeP9Y+TzzrlbkitBQndXmU4IGQPwcyztJLg6bxfMdWrnwKDIMpCfc/gcC+w9E
zIpNqDtXncuvoxJShbl84EYK+ppNOjeOlrhowLXrt8HKVdYpOvgA8Mu/ltIj/aQdD6AjdVdIW5eN
xpwPao03IMjTDAtHixLD1412HIT2+5o39EIjRrAK9VBzZ2dsHDXMQVNXbtEaO/VAqWFzIxTxhJ5O
yEM2LZHh2YnAJxnsy/PqCbaHjArte+aWFd38mskH8tODJXtI+iQ9HbcxMxG5WycKviO/+PbQy4Ll
uItGKJuqZ/Fs7hK/BBZUnvPwFtb6r1jnqDN0QbbWOk3/Q4IJstgSXOtXs0DCEe9v/sh8q+UBzfJX
S8vKFJRysJU5GSpT2jxdS9nnn09KuIJrmbT7JEsg5dyp0RSsUKoEz0qbo2ku8uLjGln2Eqr/f9i/
Dmgv++UaxiIbDayO20tluHUxl8LmjKmpw4R6CdS/MYqk45jgn0NsXEKWFr9jV5RUj6NTJ4udDyxw
qz2WH6VblOFfKbwS9i/RQ+Jpz4S1wQFqAGD2C4vRK3IyFdDdTo/armjC8kAjzC+bicGPAXCO0LwG
bS2MC3u0JlNVJCY5O4z3CRdIUQzdl7KN9K01arNlSnt3rjTX6ncJjH1E5khmdl8ReFmi5Nr2VJRM
B4l9N6hhymyCiieud1qj6hprPVcQMVkRu5rAKUvnsgb/tvPxUMshN8rbQuL6EyYMlxwsmGAiqW1w
j43QXLzlJAKoadSmXA4UT1Fbrlat4ZrW7JElsuPQD3CNEu69IMWahsBFNewdO+D3+gOHrqlaSzQI
Bwkc80Do5IiFGSaTIBzLQMKmPgAu6w+gpj9gHgUgSLMcGqFoHJqUgbuDf2S5NYFKKltcyn4L/dhu
GDLGV2QKFYFeDLSQ8UgVwJaVefwdG03X80+qJ3h/bi6Ua2PIifRrWbHkiqBAkW5XbnT4nhRigswN
hXYpgyzExMowj8l0QE3vYq97eQ7OcSM59cLDr7S4a0TQ9p+V1OsY63hH2075gZ5qQ2Ct59fwD7AI
THApSt9d5UFOyOF9+HM76VbSHhpS6PEkbj/uVsAAouZoHacWK6CfG49Ga0PUl+f8uc6KtrLiXy+N
MyZJ5Y+HxG7WrPz+W5rMT43H26gstUFrwepI25t/AXq69IStDGNYuLA4W23Tdmjgo6zrrn2woAGH
ENfxExA4H7ZbWHOFT+OfZSVUdjAJY4gnRYazMCYA/tallOiplU84cS/vYnZM3nf8gxBs2QJDnGZM
574CCLK8iJhZwR9s31aUcUKzI+LBWM29jGLYKxAkgY7xyY6XKWyqgLvDSsGhx1Z4hOP1FkG3RlvK
pjQ1yR5xORSMaN+pkRiOw+PEy1oVpiinRMSTz7T6s11M+PYFMOc30hAfVo4vAw+e/wf1nN1Y2QUB
QmLZ5laaDic0jpNmKE59x6sR0xK4PTnGlAL2XYlBIcOdG2VafALYKZgm9t9l1cVT4Aict4BPY7xB
IIK0+uYAHMKySjCNNcLtmTEtHd75Jj0NxbWzqvv1mwRFxlge67A8girInrM0Nm8cEQ4kRnUoZCXb
6P4jgGX6KNU4WMOEnPIb4gTv8kj6ojv5Lies13wSxkB1XafErjKh/p9YeULnVNnTJl5Q2xGsWzQn
77m7+mrTe8lEDvBi8U7Y7CLqNKtzpufBypUmY63ZD6TPR4s6L0KudEtQ7I/ig8QaNDWmsJr+TxFM
phBsuA1adztXxKYF/T5cYJBwgUkx702HefHy31Sf7PRHvC/0VDb3FoNNuimkReLpLedhLmTVWpI+
mSvqty1krCdlLLmbHUhLTMDQ05r61m8o2m252mviPQeBMiQGhLPxczvrW/BQUtVXEypSHaAEqPN8
89O1ynyQiW628rILYJXZB5zzzD7fqjJ4l2djoj50NkT4I6jE2Z8lTeygvH8mGk6a9DLeW0QEjnM0
JY+AWre6Mr75nQUIDhU2iqtGnMhSy3ZAPq5KZ6kCQUz4fcKN2Bp7+/Oh/ICMMrYPzG/sqKWsVS/I
b/9AjcakTXn/K+EM/T9L2kWybVDJk5BrvtlHcu3girJqCfd/zIwFg+jRct1dnIl2IdB2CDmm2TeH
i4NHYP7r3PuWuEYUkpdC5RX/053yR1UvTwkAoTkPk1kM/7CyAzo3MLvFOY1UDKyMZEHHQg1GY4ui
ZmipwIuo7Qt7v7nrq21UoTDD2udMqkHivg9cQgaKhJ2rTQBC5mau7NSGJRUr+FlYTIq1XGjipO3Q
yhEtaLpxnD+WWOXaCnRcTRjC2aJ5E1LsKXCrFbRkXl1sZWr+78Sbuv+PXNRBlHQYXKBGnY6fkdC8
XRWtiw53zlPvlu+yCCjhsiG/odxYLzU5+EvjBG1HTJqhv//Il/1iXMbIWw8eyR85ysIxap3KcTsv
yeF56slBQRXtIBjLOySE8jQTASmH6UPywt2KrdYMaBpKg96NQyJmDFAKeD4X5m0fvjnKlxn2NuYN
6AX2efArupP58PzM765siFeoCpNZapuGlrG2XgWoVdh1G8G/Z55yUD61YHW5ktdsdMHBYIhCYkiK
tCCnE6jNeokOHgtQ1FGV/FKqyCOVA5iDMbUeRDUWFtQH6gk4s091ntojW1EvPnDkaHzIASqpoLeC
SIKwL1wVzJWMYP3eUkOxScytQR5kOaQETS9aNDXwIPvMaqMX3DvKMVNHKZ1c9rB2DdnyH8kSnRGg
D38iDoTTrbWOTySuG2TYuB6HIlaCYM5siUNo14vBZ+JgNCJYA8bANUAxmzDYQANDZcG28XeV2vjU
eLadXA9QpZKOMbTPuO8P6IhFJ+fXoQML2+IerkdmpeqxGQcjLJ1ZEhrGLTESJsWG78xVGHgKfdwd
6odCq+KYALIrRHR1UJUFzDm0ShWOMxoXfkcrz0i+68BliJwjMa1vWv7Wt8iLtLrJoVbQzWsRPWRL
jyylbkQOUESYp16KKIUFojnQS8r/TGN9D5vd96+5zrZXb3TYdIsOlDRbzzAuuHVv4KLlo330eJDd
Js6oKR6Ep7/JpRK1kk29bG393lW0DkXuWTOhX6/VogamRdbxhMwTJnk9VpOXDSjuXBLsZYsKCnb4
VjoB+xb4fWczLn24RR9ea+mwi1CY4rhiSelNBT4BXILsjn/3wu9cDVLf4q3TZPhf7PICkmmZO4j5
ZMJn92Pi6PUf/fxYCd6rxiqSJgaXJFqmpbz8+IGSFwzPP1APlYsxIrcan0FZWGukPx5YFXpj+Dwx
JkUR3r9T9GVXxuH1MDjlJUqhKzUgN5fVShhCz/MzGjnucTs5JPkBJGqDOgfaAMUMFu1/aIdfwiws
WtQry8HCIbE/emtVoOg+1GWiVWKPR8BUP2QYMPzyeF1y/HMZo38tAKJWG8O58qgAhOv121PWdZ4t
/3Ymj1b8ZFJhFoMz/Xh6p+0Ubh9agoCx9SlQ3h8deOcs/YIE397CeIEIsmLjQiGV2tcaL04CCULJ
eI17aUVyNfCSlIqxaqKcpOlZ5p8gP9Jti+tFvVSkhkf8ijGAm8KmDZ6pPAOF/5rZOl2RPTJtwtbn
RJhkCqic9TV8r6ceIVc8q8Tzd6xm0N1GzpnNSFJXOmZxwOKgzF5yP5fOQ7GR3qKg/G7GUh5U03MZ
FWvxKkiOCn4eg+s55FydK+tVSY9nKQg0fFf4hl12at/vwx0tz0QRBl8Vjt4cvv//SQRVfX0DBFct
sPNMGyTuGTGjnhavgZRDEmHVYymMbOUtHpeZOhgXh9AsnePEF8h8y/KCrXLpdzDt41+Z5wgnhM9o
8KqbZYRwTaBBXBdOi+6mOrxLe860UOHg4+NQ73rjiUXuUMHUiG4pjpcnq9sHdVZbW1mgz922UT/R
Hnng8RTBWe3e6gk/r44O93BUtADyWaY7NHBpzhDuGz9gfoXOdN2eg5dkW16+XOH7rfqXQjTNGqsA
UtEs8quBsIGXZnFGlOIQYJwb+mbEUSpDhz8GBzYI1up4TjqCH2ECcmVfrmkAwiR7I7n6t62VNlFU
z5AFy+qKvfpk9QhQnuiGNxv7CC12+irZg8DEOw149RHG5jBZwQYJ/lnE2EuxUvf+unk4KwPWI67E
gvJiHpH+ypJoGtppJRoVCGiYllMHPu/OyTF6c83sOoAxguX+VDjBJXzwCvE0hWZy+HUTuXvEGAsE
8lXMb4MD3a8Nxp9LmvTdAmSnYLGl7PusDoYqAVc2zbqmjwFeNEmN1PxlVpdRPw8LVJGz/uSj4fQ1
/duzGR8XPSVTLpptrRAGFVco6preZsQDgrA1Q57yytfYc7lpSosMnrCMEi7ktot8EJ++rUHPFCRy
KH9wkz+n5FKOMmr7NWUDs4nMK28OvS+tkvaY7W0tzVW9LvE4Q1T4Ud7lQX7aUVYXtFnDSnJVBobb
wlHG6QIWYvD6RzKmIlehCFJxmhccnCsBTptC/ui7igMCoNUS9fxfmhwJiVcHxioYvYZGIOKcjnEV
g3bsTlA0hcq75eBblDyfJCYlRQ7wxsaA7CKcwIb04HknsxFRIEObAccCmJmVce3EWv6kDf587SuV
Z1KvdpT/uJLzCghmr5f74KSG5pFStTIRwy2vWPmCu6wrcH2nWTGz0vHl9n0ujbXxxDWJQGNGVKTU
RXk9K3SlWdbH+3bHrFErG5Up/85mT17ZS6aD+/ZQLBz3fiuzOVNgMjxI6cWEELU8oxS1pLcRh/GW
FqWMFu9kxITQxA1LE/yqVnZt1m/fZOf5sp+ifPEmnLb31ohyr86Ormabcp/d3rUGUueKVNv9+XoZ
JkZJB8O+Ci3x41appfbknvzss7BezOILqd1nLUfVQBs/xRVqL33Fxa6QQvkWoVzUGr3uYWh0ECGy
uP67oY87qCobSXQgjU+x9TIHiWSd+X6upRjaYdiRNUbsbsh+qucuIybXQ89pk5giN8TlNfQj4VDJ
bIL1D9U+YUDuoYngev4iPrcZzQnK7+CFpY5V/dHCjqZbuRylNzRGJFx/xzJTZq4U45yl4/9FtrHi
6F8Djq1zFWdJRRE6kqqlqwNoPI5as7T60D0HR2n5WPPMZDfwPdloXK3ZbEhbj9lBLFLGQlMqpsKx
K4IrXMqT4Nm6u9RMpyU6BADypeFCf5FbQJYwAix7qHIvYWC7X8R1mLdCgsn0dPxKZGEZF+zNd3zs
knijwL15sZoz7GMhyGusZicQBDX9J0v51QTiIvHl48sYKdXqppQSQMXPoH/8NIBHRYBMdhy9Wy64
tkuE6mjTOmhMXO4DODyltxIlAvww/d9v8Rie542eduxt3+my42CuR7IGpOiLvaflbGmt79/7NRNl
xDLfPF43OLqE8QhAaSbtUOIr7eVvuptPBnGpWICy63dz+IkwZg55H+kbumKvqCDq5CK3ltIgY/pg
u1jd0y84q+CGcm5dnfOoN7frEKBuZNW++Ci1dFkJsES7KxmMhAd4xMsADZy++HgbpqD33MTWu/MW
RcdfckEEBoNq2GCbd/mofiP9CBxnaUn6vcB8aJJbgCJUzx437UCbHzyhFBssjsm1EJB9aooFI/aR
Bp48Fyibw2y51has/8WoBvrwbEjKg8SUdZUlpQZgCC9g/99k4tHX2MMOUQ6ldnmGtui4mT/W0gDC
USqssSM9B1P3D2hnCZ1+AVqdRfcPHjEyoyM4P+1TMgOc95vCa2SlEVEU0K0yprt7xIwO+eKAPwVJ
FOXxyRUEx6UTIIsa7dkQcgIUChf0eJaV1GFWRazYHVSDRrpknRjsCI2bRimskoz5lBtnm2i42sUS
pkL2qBMVoinh+sPbnJBHRv23JctXMvLM49IA84YFwo8x+w9+pyVMGldU+u5RaTdOdd2nE4+QmdFg
VwmAVkthGroHLmQ0qq+jtCRjOckQIwdpBqRJ7GTzn+7u3etjj8JiIpyu0hGKQ+WDSs0Gh8YDUnr0
Riah68jP8XYpVj/kCWIvriap8sga6EdtF7ImZ8mBuwHK73Xga36D7wHuArZErzOquMgsXf+bJ7wC
lAXnBGhuJsHgo+4Td+FTgDGZrVjxT9wNhU7G6aMMHhCDnC1awiqs1qvZnK/F7es6nYIPvKPC2hE4
a+K1qAXVhkVAPNHYj2CQrknFVhTkdtgSinW0jX/wLDj5lPKWlwh85BAMZObfoOpB+AwDAcOBDF6D
LSKk/cSmECde4fuMfxp9OvQoPW/0BZg+bZK7cOhgn13FPS2QJ7FsQ6aCv9BMezobXxzd86ouvtOt
UtGXVUmAfnNHq/tRvrEJRCRCnB2H1SeTEe9hdbV5gBzlvVWlLwck/fi98GWLDIuRym6GssevDA/l
/sW+rMV82icJARdvbgh4zNHVbuwP7uIaV5gCtfBTU9nzzGfixNj7X7QkSI+YTz+QBg8L0DsUV7yG
aNWQMLFhfA8/BfLQXQeiYuhcAaxQzLNEOMeSCAcfH/FaL4qp2DtPcn7iGU1nr5CKA5hM+GJD+D/q
QSzuFDpkms9d7AA55QBcWK/WwjxOHfVNXWA9q1OfFhYV0zgngaFsdTqTCkuZfkgha4pQU9OSzWxN
M1IAKtAX7Po4F3YyLC14pN8W+97FGu75Fo4PkvOGKaUPQml3JpHswaO8F1SGCwbYJYEOSCxfQV6s
1U5rt6kyCGOPs5vCMf40xS/rkN1+4td5qLosIXiJV5ScTopb0+pAWbzC+PE+6AxzT7PeKGEF6MhR
th3GZe3mp16IpOYg4wC1oLwpu58Vw3C3Kv/0h6OpOFRBmaJNaK+J9PBY13K6+TkeHGCPXMLjfhIf
vZjFQaAg+0HJzs1gd75wkVIqfFGwr2zrLQtV2QMx0YcbM+hMzbqOPUyQlspCTdcE2H1xjfKKCuMb
xjMf4PdgLj0ZVtOtK6VMMjwTCrpeY3dFRlXqtjcFkjkQSYxAdH9e5vgdq6YOyPw/IgB873+ixWwF
4vkk5iYbcum4Y04VEeALu5EEU+CVcM8bA74HAiuYPzkk2pWRErfUs8nIEpRN+QuXas8miSGuAobf
r550tdKYV8S408Oj3DLdU4+u1IxRS6TIWpSIJaJ41fODC6zMIajVz6Uv9O4L7OLS8a4FZuwf9S9q
Wyw9zgO3MaFNyiwEV7u7sgBnWjD0SS6t/0qCLQqnE1ChMcBb4szpVTjMpRxHANYA7dSr1j9VX67C
D+gUxnxxLNhnlmvOv9G519bIVXv1K2Vi+vDUaHuFagySkhRYyCneEyjVe/vnLaG/ttt5OsCNzTJm
iC8yRKokquIYOHn1cR705GgwQ+zfKJvubo6oMqNI6vafT6cbY47kwMEkTaA6J9PkigpQUKLj94jD
PcM0cZikVCC1ubkCwyqvo7G6dbZslYr0EfFMqr9yVcSuvyXVj++d8srRYMz1I5RtyT89Zp5zqWGC
EnhYKh4hcTsvIdEg6Q1UjVw1ePgLURyIh6kjDnvvFZYEEfYpeEmxrD71ARNMQanwCYg4Iqe7An+g
7i6iwUrfa81FO8fOYiDkkM8PkCCIpJY/fX+7S1LykZjgTOTFYCde7xgTN+kvMcRL94eG4QPE1A23
HcbfT5olgQ8Jyc/W200IYN3FOXlNGP+MZPLIFnSY3czyBDMJZt+yLJQiBGetNTG5Da55HO1yAx6o
MZGz/TXxzA9fdS5Zzwn7BwbolNrDSJWLf8g/Uv4GS8JAD5/gF0ZrvJy1OJnMycvtQsx1hIi6YTpl
NzqWZMSBNnPBWyRZCbz/FWijxxe0D9DPlnzw3jydUeXyWIc5Sc/ek6duYIgUEkZH8hghORsBHY/e
SrdE9UM7Ox9wYFfOKq9XWT3762jRz87K8pBTPZYf4PQbfjIMo6Qoc3l1G16Jk3oujY9w9ukcW5HJ
L/b7zELWr1Wa3d1Ntf9P3INhQmWpTEGzskD5HvnbWF5ysdBFcADiRCMDngGDMKbcMkIs1ckE4dB7
MFUOADS8WGKQQWpVoXAgcNGxjX8czhIX+w7jHZ/AsRJSaICNpKKNnrSB9C24U8k0bfaTqF/2ZHSW
qIBHVkknzkg9Ysn7Eynba09xki2lzvg/pIosAioYNZowLYJ7uZNYuGmdiPa55XqfzvFWQL0+KSOu
eSTyK0BtuQMq7FqF43LJRpon3g1p2/kCGC1X11BEBQDxwotavyqW3pT8q547uL4iDW/37QAJ/WkV
1eV2fVPTpVXa3S9FdMjgcPxYUJqjQ9JyPHKx/K0FkjubEcCHKfPL7DpkWszThUbkbxuHTGcF95MQ
O0lFJVOSJANHpx2BIC3TZbqkB028ZCLYgMZo9kuM9OyGCaqQf8X13ZnK1GC2/ini48sVQK7oSGY2
UTz58LZ1/FEgCxVN1U3+l1hXfBmpyAPYoMDqjwewekADOo27ExT//fKpoS1r6yyCzJFwrD6Ma6wH
oNRjzKC6vUvQMMIzD4Q1j+075nYdn2Lz6f9U7Y8b9G1u96PKIx+779unoAV6Yex9hlcXGJZu2hsk
wAsWt+scOS95jgU4khUGsL9BpEgnjvQCErR9suejgW2y0vERJ5/kH59+hKWodNsREigXbAWHZe/Z
sa7rgBBiEXVZkVa95I1OieyUoaPQ7o++baLvGqzmd+diMmvByMzWDz/v6ttz61yoXV9VjnL9jXuO
ftg2Sm+CmaEk2VpVa0hZfaDeWhVBnURi/v7hUlrbliHzWhejDpf4X65xQ37eWmoKNYoPXy7hJoXY
6QHOVxN1k1gYOuDnnsoE6cnnhC+tqR5hLCXiqATfL60JLGCDRl9f5iYWh7hlzWAqTB0NSjEVvipe
RUAtYilZPHublYxqfP89c/j1yOlm6uUPg1/jtHl6pkOqcb29JIoKRw9SeBujD5loRQc/KleCeXu/
2tsXi2ZtM5Bnq6jJthfad8PtHsqbeDyFADKOcL42tKqV1JzW0cNs+YJYnE9L6pwamv3gz4EzZ0Iv
9+UYs6Ntkw3fNBk2teiBqXlrIxc87ZNx3RNFZSZv0kGHoe+PZ7nKCSqHLXu9qy4DJEdskDmG0zdO
M+4GHkkeipPhyRU8xO3HyHx52E0UzpjdcDolG2eKrzaItlOmDOtUGZVRYgUnJYhmeKDWpHai/ypm
MthYx7dpr7ZpOvJBjIk83TC3YfDtZamb9i5vZm5++ic8a/V7lRkrfOwn8LErFv9wU/A1W5rFekfL
aC8iWzPXJZARjT40r5ISI4FMb63etWmIGvRMOC/2ZBV/XcZPO/3NKSUty4Ch3IgPNVJHsijfhc3L
G6RZlav/nLIlklujH9iWv+mkddHzHHqd0K7Bu4u3h04n6Te0rBIlj4nEVItpA9yorFHUko9t33T6
1btdhf6hRy4CQiSFuMYJmXQQRxPeJ4prBHPIlCJhC7aHPruYp4RXplNJvarC5kZQpJmqZOSRRucg
653RlUIwdOswf7muRsO/9RzjE8Uq3GtSr28+vH5OuWtRI8jyq57t94M//E7ye0buw7p1ogv63xPt
biP8MDe8ZQFXQ/MsF8g8LN7sFHOHdjFVfeWnz0d/f4s+63wd71s4Sd0UHX7zVIFsY0+tBBhhFNtc
3osFt5SS72be4be8qNbdLT1OtsznnNXp4eug8uW5JppqM2yDMIgXcbSBdMXuZw4BXAjrMWcpLnm/
y0fSJTn14w/stHLA7HXaDyxtsqVAnFasYCPjfrg5M9EpGTAYh/tZbh+273n1Q5d5c97mV1SmUPFQ
f9E0NSq1d/EDTWqAmIsnYV9YpZ+X9Y7ck7J5weXhkfJ8VbF6SwsLHLvkxLC2hW2duxQYbdRP75cX
X2J3NISP4WLhyiTlzU/Dg84SndlQwylO0fxHmw3N+mUvmqK1+1ATSIBolNbGnFar+mY+HWfZhhDk
tbhrKNS6xbilboOmtE2cuV14B5L9msYb8BSuKLlRUvVRak6T3CP/QRLtf3OTnfDHJnRmggd2xstM
Z5RgUCJjypFrTT4SwzP723Pg50n5duvF03hQ2YBgTvRGQZ9R+qePl6UNcte2pOZIMmJZRVpLJd5s
GPYEuXEEDQ1cD3t3dXAlu65IHm06c1mQkJicJd1HGA5F7Tz5jzy0MBp3teoaJ5uGvcfrDwMJhQ2w
j3R1Gn9JJ9dOFlvmr9RrpWTel1A2YRcQFDMVAwEB9vD2B3mulq27JMZmM4rwHNsLn7mnynFsoopL
UWaQXQqQi8MkCfymk3CwAgaX9jWy+t7tlaNOV2YG7YoSMlEygzfyWbDVqpoCA9MqovqzzB0FZJNk
nwvdIgoWZ7c14336JrA5A1Z/188rx5lIPD0v5RwOIwwZdDcOW/arBT2yHyxsFnb4w2heVWe1JOHv
RQ6wtJjCVV2uvZgLlJJjVodLocTvgt+7p41JQRHJcjAUYKg2AwzDrug6RozJ2YRJQYRVHHGOaQXD
QHiaP7sI7xkYY5JncIew6OR7wPDPzVoYZWs29a/ck8SZSUMc8uLD+suufCvgfN5QkHAjPeHIngr5
8UkRtPbBOOZt4Mi9H9Dq1pSpVxDxzYyMIXlu+lf+XnXqXmD8E9/e8SROxs9oKTL/RNZFm8AZoBgP
yoa6vAWnUNNBXIFP2rtdlpOxpaipdHR2m0TOdqWH+66ljPL42jl+/NK7W5dGfu1Ai6nL0NwjU+HM
GIGe/vgphH3DL01aAB6VtI7Q/Sr1UnV3isLF2zFluu8MvhyyOks51WYyPlVu6XJk81FtWn7tWSek
B9GQVT1Qp67UoC2huctjsAK9hWgSSSKT73SCgIcCHZAdl2zFwzlUAAOg0tyL6BfD1s3pkC008LN4
YQFy9OiB3GiAjo6Qmd22JC/lpA9+uRAg7Li3oi5377XMRAQXYZau/fbIEb//bHEgcM0GM5+9Awzi
T81Z5YKfTcdJuJLvv0U4snHGQhOgkb9jYrBSqr9btMUwyMf2nU064nXYWPnhY6gOxQgX2nhSDwkh
dz4obACvvGWbM2knT/2LjI7E8CCWlzKaBSNI/5Px34pxdCfHn4wwm8Pqqx0UcYqIIYkx2HMYwnlL
JCoCEy3KAx1bqQc8ELoGphd6mKdZhorN4Nb8KoD0jX+rpNifbsSsdrLAAOLambv76VYi4eEiDEgl
2sIOYI/op79fI6rg2Efz5Nmb5stNMQbKjTG70to4eTmCnwQ2MUraq4riUTElpi2ET/ddO+w3bQed
yCPtuFJ47Ycqr1fuaLnQYwXvwJnlWUKVm7D2o+Lr2w2F6IdllKVWqBnsdvzhJxTpxVvLdLgpUHeL
bDIIsBL7sXzqUE/XQtmSOB0amL0eZpEXGPXk9G0+h+Vvm6GFPN4T0Ci8MaifMC9UljmN37dK3H0/
zpWTx0aYTVHEPL3+FzSDOaMZ04ck8nhSmzjz1oaw435CYTHDhhWEU5+6qRtPDIZC1t2OmzMdF+yX
nqVLZXphrEP9zzqbXFzt3o2ioNcrnyNL2yvDGwclnS1I1lNartyqe57yRTITVGWqdgvWJ3Eeeww7
3T2gqfA+HW8HZbxJQmHtOgNno7VQranZnnlMvkNa+N5p2FmM6+0PSQp2cn6YH9kfkybZs7JmmQFo
3tDIBHmV0Bzw1FLTDMkQcFpegZ5IoDiz87hp4iAQJVwe43EocytxTcHPRym2SgbHicr3lUbjQ8Kv
Cmzm4wmodezDnG4r9HudOijWGyQ4mQ+oTLDNuqb/FvUahU9ZgMqoKfouL+iStG5QsnTERq1HWg2+
Pu+z1PekO+5Jzwa4UOgAY81P8tFgnlvuLBvo1Rx+WIY1amHh6onmmWujIA5MOyeSP1whx987mGSe
HmhZtDs99IxbAXdydcgzAA7axI+2UCtQf+FLUgiifSKRPxmkf+G6eKKRflYvv4k18zSCwDjyLhpC
yxj+h4bX1A7AzP1Zrjp4jv0aVz/vUR0OEWfC+K0q0WUdZzcgJoIOe40YQOeMriEXY+JC/9smRW1k
ZJUXE0Cbd/TLoq2eAgCFlMOaTMH3DWPManRQMfmjlJoogsBOVFmgzlLIrwL1GtfLhzVs8OvqwDAS
kmI+PeMo/s2gsU7J08MXr+IROQmCIEDwemvk9Us37h04fkQbq7YK/++KnySsdL8l0DcsgbmAu6qQ
gXuavc/eb2XqVuAoZAG6+XqfXGe9bkLzxH5kYC0e9kwpR1X+ByNjtfYajjw4pUsktRxZmGhDFOFx
KGscqA21U2I8L14JUpf8FeCGXwmJK7Yfr4Bl4IcwzLWuoJjHVJDgdNCRMwUZ4mWTtcRWjeCAaIlO
5WbL7qmktrFL7FdLfzclaz2lJaacpMSIb+hD9X381q0C0FkSA+qKiuSNgCQdmNFI7u0ufc65DWBE
TqdDaZTcywOHmUHzy6jnkO1MBRtszdH9+lhLgO3QiFgi6GFvplniy4fsX6vc242QjE2lRjFhvDCX
HBA4R0JTCmgNrVNibt1Px3BrONJm6uhis+zQWOrxfjzU0ddgDmtmoerQ/ggJakpQsJvdzTzOtsi6
alzrxcCkf441AwXXl2m7PeKcIkzjHJ9IfbYdR2uQgNhaqZYZ81NWHqD0j4+P+lqByL5K4Iwy2Sy2
tBKOiikPIlqB5hViwtRsKHVK9LAwH9YucsaPnlWXo3/g34SlHWrD0vI6Q9pAuTAbpfBqmbfQLlC1
Lsk8jWHBRxUNg9+lk334AgJwaljVqRG0yMtaPowHTNttklJ0A6uQN+8CH4MVEf2t3dSk3LH71VCI
J/fyZT6OJ3PDJaCvlG1LXwCYnw/s7ewKOO0vX1/tobJm6A0E0RKA9KZ7Tbgr5BNkVth4XT3tTjYp
2uohSrBQawfuxU9yHRjU9GdbBgL7Hv+MF26A16e7UACUIkAIBPKIFpePkfQCs+RwVw544qwvKZjO
6Jwjta01euCh67o1CaclNEDZbdxmf4QIBzHfdbiwBHOW6nK7rAZ1BeHNvf9mVKUw6RYquiKokX/S
R0yguyWYrptocM389+U4Od5z1Gpt5yl9CBff+R5xvJn/Yar8yeLLw3cGQ4sBMujwsfnyO3z+O4MD
0z2RaB6S2XECTWkRR+W0ARhIZ2FaC+Rm/I2kM+Wx+GsMOuDcH1NuFQc0BMlULgaEBEGR9Yo/G2jc
HmWCtTBVVs3hRHfvRuJ17tkH9RLpEBtTdoAc/ceYUtD+1Ib5rprV/Mard3ZRiE4CVb6BJGrjOPS2
G6cfNc9nHLKY4P+KHOK/9Sququ0eJTXR9BERk3nZgIOG0/rwpgG8cII7tunxAQljgTZXaApc3BmJ
SjMjhBWHpsdzx2GgTJRDY9ZKZ8UoVJQWi85Z8yFl/oLnPv0SOHc4ft7F+tWA9Mmzk4FQGbH0e06D
+b06z1+fDlhwJsESqHA21d7yQ/0SAj2lFiwqkj3jWkptxDgSFTPb8q0XQ5IQFARNpEu8P9PgT5Qb
zei0vMF1esSLU3xBw3JtLWpbsoJwvu3tN9GnaMyKtHRBL+87JmkD0zb7JXY5lRA1GMvYuMzKRGjt
DNmk2T5RhcAGmq00Q75gSmNTGpsDK3HGvNw7hsW0h8KXL3XurZx9rJoOn/ipsS1kvjIniQGTia7c
PXLbTMWLln6k1P8AjZ13aPfb8f2USSrv+a1kZvHLrA/8BcFrE9/1fQT2XE/yoetkdgI9Ud1EF1/E
SX/9d0ie+tOyiJM2Ly50SDOasXVEtWRdXpy7XDt0J3UL5UcAWHfSDTE/rtCFwkXSWYz1IonUn3Cg
pVY7IzXAybJgNAGlqJfaX+R9+cWaylx2ynnNe4BqLs26kJ1N/K/J57f1WzBdU1iv70UyQJUJ1eSL
xIRbsZgkPbcJO910iCyeec/Muhb9L0TVbxEGfwD10+OeR6BEwwW/b81MzzYe/eRzuBBTDoiHeU+w
/or0vMP2ZFHFnLbbP5aVsIYGp4UwNs/nGpmN/QsFj+e6Ka7N5vdGwwq7U4k/nYsh6IGbHnD+9gwb
lSLLIQlQJvu4wZ49aj4xUQ13UoTtwnMeI+I37zYaaPJGUe+PsT6w011FBemflgSu56o31uCqFKIb
g/VJVhUQ2VvnfeZzTke1Q07YZ9hXdgidlp/NzAAC1aQSEhPyI3uvEaXu/Mve7lkCWapM0ESWY5qb
/q4IETsQG2uD89evr0QzdkayMpdRi1EHidct9UvDw/Rywl4vhH7HWYHCXOq4XpTZn8h2MYZgDW0H
3se7Yn+W5Hx7Mohv0fVDb8Ziz9nRN0hyMIIAcYeQZAP9rt9Bbc7e1su6tW1o46Ig95ABK3p9+GIq
QHgzp6UBhJstqYNxHREXWjQcn6i6ggj9VEs9qSWsKMYPr1knth1L0YtP1/uFyroZjUMXxDhObuEc
bBg81rD3wE9XW7hPK0fTr9tsAT2j9O1xni4ozaWOOCu9LHXbQcJD0uzMpPITB+IUey8EBITN+Tct
IHq7qzsLvxzRX8ZzH3ffOL+C69bOSFLENHMzWWrwMO/2QdoSS540OTwDHm7GgiJQKsEdSrKA4BjW
lWAf3HgfmcNCWjEpjW4/3BbTYXY/NKDpdurcIXLTu3PhTuCPsCENn0JIGJsWIegappYeR3ZwAlGG
fObO9ssqvt9ry2if2ybVHF7fq7FqhsSUKM3fCbuxK+gJ5LsRNK2f4mkBKMmyxZyaBFuP4jW2yqvc
53JFVUZEsP8SaaOhCBU2tTnl6/ueCmzWTfwZCVNZu5zBNNC+s4Ysxm3a+XVYN+kVW02+vHRAlncm
IUEm+vqSf9mlQsVZvfSYwVnHHHm6xMlODuOqULbtIbYKiXoKjgkLQCa5kBpqIMCrPvpMAxw92ODi
BpAXAXW8GT8wytXaPVnbCHg5ddep1WBlPkzoV72+xSNMQSZK8Q4QUbpg1/RZoi1oo+mBQJGAh54v
bHEViL1CF/BlKn/X0thexEDHrP6GZCPTFI5I5u8/UqLkYTNhR/Q08EdNW71GYQ/LhQkRMVrGt1xG
dreA190kPMMMLB/+RH5LPiex4Hqx9BH5168aOkchdnlWIcd7auublF1ytvXhV1SMKGr2ZcoHUFsO
fkdqBcbmgC0KwkUjP3yoOO9Z182fqZsSdnyhvnbpy853GZehtOO2H0V/WyANFDYK+CZ4KYRP/HpB
ZlqpnKXYBjdBhOoxRfRLZrC+JqPAcwXcFMorDTVCBMvKq7Pm1Nk8uHRG0TlnLvDx+seAB9Jn4Zxb
hX/KPtq3o2Pz8s5XzkfrJGkP5SFZu1QXVLGwHa2lu9J+I7ylizpwF7a+Pacrz/Hxf84swLLNEGEQ
8+U9ZiBGC4HLXJEWgNouQe+bahccLeZeNs/1LXbYPm0NaUBPknWWSMMj4qGxcxH9a7g5owJTKjtq
5eMhc33B3x/07E8+p8wKnwRWYLwIkJvNhQ3ZecUvQ3tXWabZ3y1Y7EaBrCaWQvKSlzNNnFmBLWmY
tKKHRsyrmtFr59Obak8sG0jQwBjKdLB+igxJqMB3g5IOGay9dLp3564c9s0UDQq8ctxMY1abTrA1
2uKdjHHSruLT6i8fwgY+/LAL4MlUFoLr1k2NMf36iQN83SPn5nXhr90sESsCOoaSctdhXhY2R52R
iQoMkXfVV25LG21Tbg3CQgxck6XJpUZHxjNT7GMZlFu10TWTyBoeSMcEtuOloC9K7CVO+IfBYK3J
53z2IG6xNzXNQocdxbaRLWaYQmF56P6Eg9dEVkNpoVc1EKhHY6JCZ0XrM0oV40sC3gItnJR+zb18
2kd/eWQi/NPwX/euNVXYS4nwBFR830aKokhtQD4P6JH9TXP/v6aX5o5HcrqYDJXnOyjQ5o0QRAQB
/QkzOBi31dnFDxxiFWeqPFSKa9zvmiKpEDk8v/dL4v1UyyOcORFvfnGrJZhIulgR8Hz+3YQtCzmW
fT/S0lH83PKVy/RXV25rbaVg8HoTBVlFa82t3aqOcrsbkTUWku7qfrQZRyoM3S2KQVkkKv7ALcI4
jn1fQTtA0v4AnbQJ82Pqb1mmv4U1S22V2FkE1kMsS0l1k4Hl3lKVq32tEOyULHQ07XIbIBp119Kz
K68bt3OXdOn7Sr0/OHMf0nOq1aF02w3CbA6IHu5Q0ykAzjd8A7LRPCY6HmtVMFp8lDHYwIG+ppFU
mAAK92jrbjRuyj3Drm4ra3wCYf6jg0xymMYTUn1edXq+j+X+78tFKAuBEGRRaTJexwmF9clkndi3
uXguMrepdnWUmWatZY82SThUxQml+kY3UFZr7ThWQJA9YhOFyIT9edDIWd4feOfCoHeP5H2pWv8l
6w8KOLy7N4JxSz4GV5NpAPrw+UID/f3Eu6JPH3GP8NPms5ZNvH3o72NK9Uf6undtQrR3xrI5t7C/
5uC7mUmY68MypMdSarzH+saiSlMH9wLFQ5ixxoSl3zAIqDbx+Jcdk7W/8BQHkZOsRY12+oq7usDB
ucjFJfsjT1RxDH9utqge4tcdVDja3nL+VmY36UK/j/I4n4nuBdU5gttFfB0TCyyK+cqRZwXIbVx3
ih0zpN5GzM3pJi4PPYJP0U8cu55moXVPeVxrvRr2wi0HOGkhr2qrRjpRPeiknFJwUe8pDvlWS9Ik
VvO+JNWBX4rQ5GsoImWsz8rFWG+Zo99UaqyA6PJkDGKpIuF3N+jX4JdODCi2B1UZ8gGZMUZKIMpy
1zmaTcaraKzOijQj4tH/XUs/6w5gbkYZSF1zOWhQdDLzzx71sdNITuDqszx1JwcxME69d05F1akC
2Hpnxxm+IPA8+Fv1WS5t11JeVtpDgyqsaMQ70BS2u1K/Ekibsn0ZYqqWWXv3g5nH5W299QUu6gzU
qPyDUsBMdKWtva4HpoPfat7VG3FDd6uHHW395/wBaShT3vPNr/IY0P6MhqvdZvJC9KIlJcl+/P0t
2tKYm2CERCYdJWHv5YOsRJ8SwebDr23FvbvSncXOnnFiKQxYt7KgHIPAEB80Kg4U/y4WlC/6D02P
vBAu99FuWGlaxGF9PdWOzUaJqhVr6sBm2fN/6SYV8uXkBT0ZQA0+BBm5nyXEFzXDr4PXqLe1Apl5
cJZ9Yon4ZUVnn2P8be3LbT+AWgHn47CFe5M41Utc7uxLFke4Jei1iWbl2wIyERTedNZLFjCUAbfd
Xt9gVcRjGyQCNnHQlTEUTRx1PPDM23wW40RI34BfunPoAGq6Htnm+AHiQUX5TVGzK9iMjzc+D+pv
27r5x/PD6ca+jMpSjhqeDMPjBmXjFJild6oYK5FmRbVRSZrhbNcsU7rMI7lTrVIFmcKkVP5IMzC9
YUxkMt0e/HDXZ3a8ec7yYCs7KGKsBG8K7FtZQvK/oJI57r9qfv9KyBe5aHIoV8vvpMXkcm+riXBG
9sIXUC2KcQivffjUhlKbuSvYp0JGfV43zXOwg9mSgLNWgplbANEr62P0GQjrJPP7ESL9j3E/IfE8
a42Eo9QaUJcJ6eEWN7VCHXFyPFpBhDtbjnaDPKZ+XJpYVaBkxaNgiSBkI3CJCMqTH+Jy7Z34hDUS
XTwe8ClvPjN5YWkYnK7r4yU37Ked7W6+lq+iiLB+Fl/puBsg6lh3bO9WUmNkcwcuK/O/IIh5Hpmp
Hqjyx6JkRHfhg9l/OjRvmH2MxeTZ5Fjk9uiPpxB50T7zVlyvaBwgLh0BLEk1LbgXyKUfq6hbgAyi
5Le+Ak4xMKXuqBZzH0N7wYqW+vzYraVhDQ0UwcG5eOmw4DuDkoJN6Ja5JiqqS56MU99PvQFWCSXn
KjAbfVORIp5GfWLTcZep2BA2pGWtm+4pyODdWc1AxeoQmtb6IrLbVPpITMC/DnqoDa4NjrK9ImjW
4eCXk+Vfmimrp0M2zJi3V7rn5IQi1xzgVCoYsu5CAZKZbVzRNc6zdT9OC93CvGK0KKD7KTJrdRHd
j8xt4AwuW+759PUo2eJGv2yWjyiP+AhOLSMfoJud/BKNhnRBKSvB/98b9FP0hTflu5+TO2sbGxXi
TQOp8jBHgTJ4h/um/5i5fUgLv6QQx1hd6/m+Iti/nEdFbpR9FQuHK0TK0TLBBuRAtVWNs+zOya2F
yDkessMubhzroRJ5MyKSQTcalGPj8QJwjo3G0ZnBtOW57bTtY0nMchxCAfWrnas+ih5RU7sTxCX1
TWbEbOG1nFUDWPorlQzZ88euhv2rvDJ4HE0fesOkJ1qHBSRG/kdn8/pRmjA7NlpJsVX8O4mRzdpJ
K19V/mxMWxuth0zuaYYg/g0qjJytQ4sUuOddzxqe8c+Jp2ZrXE/DHLb1jPB0Dw1cMCQkHSl2buRl
13/FxROCLdTMWUM9H0aDhF4EY6tvn/2hH9QQO8nIzI1pFvMU6W0EV6drP/8juWq4UqS2ee4IqCaq
qXlGaMgubPG7JQXjyyhYvZdYIU+iIj4d5CwgamcoCdYYDS5M2hIAGXAGYxUq5mq81huQfcCVcE5R
y4B5slhy8FsoK2hTCQmzLax/1VvPFN8pN17PJ9dy28RVVcZBUV9fhdPLkhfgiBor82E9xNE7ty+E
+8dAD61yUIyK48OpdQB//2JJPNdtS4Tg9cgKlpPYbndH+ez2QmRu4miHtCJ3e5RJQ8wugPOMFGlm
52BePN6RV7x/VvsDkrNmI6Lsw6VEeigmpu1GOfsae7lr+xsSZqnF6kYkdccn1ABOonkFezPwKIYs
49USw4xwUp3yLu+4F3GDdzY5plMc5ZNWgs9nNYF9OEivnE1YmPYhHTHW0JTH741yOOrZacYgq9sM
FXtK/ZH6sfcxgjT984RSOxD+8yAM4+LNo+EKyGgLz+yomKZQW36nKkvhJNtn5yCFv0Nv81PbBN5G
jLaJwtqM8a356jrUlAnNwprX4eaNpLAF+jKm+3TX/lLJwjQm5PrWmqnULiyOPcP58eRdoAYUI7il
OSuzpJWzZ73mZHSJ8Sz7kYO2Z/SN1UFhN8X5NiDe/U70ug5vX+L0irYQNU85CpaKOsKWMnBvPT77
lz5YMPWlipYlvtJcKrFsKWvJEePrYzkaW5Bhp9kwGXEaUD0O9Qlq+npaBt9CAHH21zZewzDG6k7d
Sxa0o5Z5sL/JqDkbebesb7l4/+2jN+ii7Ja4StOpfFlRhEgbHRcGOJowrG16vgUGFshfu2nxJ5+/
wkTW8Nt8Ljv9KuK8o/PUXMSlxWtoQnsQLS6S0q5LiolzY/wemYi1/PrNQd76PE6ktzuvx2Wt+emI
n3a/mwJCmPiVQrtbYJWi7KNa0tvm7QQEh04HZ3D/eANrlo1XArLOKJM00WUwZMj8F3SDGgciF7Hj
WLIH3slZBpBk4+VcXzul5EsoeP0PQOKUQ9binLZ4zQvxz7QfgMTtx79GP1ouSFyk/m7tlKGwnfym
nSORoYqlt+HZOh8TjXjIjD/K6VgLGWKE34N8u808vRudglJ399zklvQk7/fLlY1QcSo57d9L1nTI
7PILwcDgTqCnc7ztQJAjGdaHVLwgUp49QyRhX0OEX0l0bp7XY6Vcw09ZAdOfJN5AocyOzetfvkQW
OuqtBN64vB7k8FDzhpEDMXibvyYVN9If2Syc21XqSG15E6DDxIVn4YDyvWwC+mzdEK0DeHXo+Ckd
y8p08R1J2z2pytXfkXB39vhPTXbtzwOzFz7OdLfSFlNHHAqUVBdDIIb0qUvs9IosZw8GHSZsEZYP
WnBZUkZMt7XjYhJYqgWqJpdi1VnYv7MI9gAcv51Q+xPbhsd2QvNe5kINbEh3Ja94tw/ghzrIwDEa
n7b68WNUOK82D7aGL9ourDAdHKDZoDQ+gW8fIxidWaeHdCv6+3/txXsBBKfrpCshEZUYTijntRAv
PsVnFI77bi0gXqwAmMVrQV9L1mGP0vu4v79WjOi1jeJtyiozqMZ4tmaZRXRV7UNk4geZwKzrcFQv
qHbnjTPhqVibwhQO7WIf+kgHJjsr6YP+8rM4hQuiBvfgfay8oI5XNDsW52uZLDCRk4edtvB+8w8k
ygaLA57ztkiqHvPFzMfq5gUER+0ML1XJV1VdvCNe26A9oeCdJmUrOV9TFQQT9bXmaeLku81VQYq4
fj1nlGnA1rupLUlAvVGJtYhPx09gmHCF7WGvoqSzXj9c4UbJsHZKXTrWez78X56MhAzqR4M7u3OR
0J+0hfhYignTYraHT3MjCRHY14JNgZMpzUwVD+wvNdwpECXkuAwkdzBywWrtirFpho/CdpUayD+1
evEjgLTgSQkkfJ1msCIngFLNShEi+gHAutIGNrkRnrcD8tu9vBiYTtmIpiau2O0da0Eu0GmupKyY
sLOvbTYYP85nGf+TwIFM5AooG475QlA6gdochcTuo7I4lJww01a+zBUvh9aa3w1/7D1fJAuA6iH0
Vqesn/EJlhkPTPxMGMcENCtMA0k/n8VpVy0hBIXqJl7jK4O/E13G7EZ2hCoqU8z6dux4fGuXq1yE
B3CZ3MKHxyZ6J2eldmYx9xQTSq+Vtf43RqfW4tYEJlzXOIaFsW4kTNIOB3Jx/6XcGf9XOgqLRI6Q
6JNaRA87RzTGt1yADi+t8PhC+UXHwyp9xNnpSKeVwvksQJdUD9sPK5KHcPlQeEIwK5pXCXiLLCSW
kDckjP4/2fa8BtxLZklztD0Fk/afImozelGCwesWwhQ9IwVllBmar7N2h+1IeMdc+ajDOWdrkOIw
V7uWZCwnD3q3QSNeHJalgfgZKGWZvk50S7UE2vIjDtF2P9Af5sJWh6a8WKRySwe4BrC7HcjvFD2x
LUSqWGBu+Z2e5npQHfbAqFyoKjpfD1xDHjUiKn4nugr1dGIjHd0RbHN3VjxcSpheC8nslxfbnj0s
m6iaKXJEQ3etFGStMria6IuEL5w1pqB9v4KPsPCi8yKsJaCDU09gshAOJqjtG557EnNcEFxrvbqX
qje5GtOcobE0LTmU9pW5LQodfRO0gby72/fdSgP8zeaWIMabrGs63kPx/mYdbZ7u2NaadILq1bLP
EPMaIQwZp9vkRZCMab4QcGOgbg1ymUd3MJqaQ7d2xjtu7fvy9gdOVEWS2bUAwR8sLsOBW53+dP7O
9Af6xj+/7C2K2KggOU7FVti4Z+HGzc4BTBoU1aIIc8/rvQeHQxRVz1JfB1weJVaDzdc8xxZHdIcR
EtAwDrpEENYC7pWZDytS4kAnY9crjMXzAByzkx8mH7SrinzvSyBdT6ISyTkO3IA5IfSsEofl4vgs
OPYbWhwL9Cdznqd8yr7xt7AYSVn0IZWaQnM8smitTHrF32Xim2vUZ5iymZO7T0AbiX9vTUP+CEQB
JcQSm/YFz1GT9ErgIozNz87W/1Tul49PFwjMuXFaO7rP3S1IjDui55GRZ859lc8sE8naR2bn+6NC
P/ubtmfGu2xTRXijjcOhXmxj4KxPC21PBAsI7V2TINoNSFvBXgn5tBO1HQYLGJnrIfS8pCbFwQ5B
Yc3E/FQ//WeNUQo08hHtVyUErA28Wqa04W1K9M1EI+CZExzSiWsdA2BzM+WedP0K3ofQY97N06Du
U0TijNgmTGrDmqVq6BKhEhaZyGpnkEP9Qm26PHo/Rfk58zcsv+3Qb+LaiwCC1gtrFPX9d/mecK51
HsrGAx8maCKijviOdEIKwTolA7RIu3ofAOTw4CCEEQmirwt8VpMxAqwZahXHPSF409DidfEZ5Zq/
Uj2ZnK0W5hNe5L9ewf4e8LGg7PnMhcpQHKMikQfQd/Jm9Y9IJVDK8DL7WA3mRqARGOEOLLqOZ3PG
sqoFWZFSHAqQ7WcuZPaaywtuNXycP2/7uaNlKk/B+oa/djFRk1Lfxi31URnCXX3RgNjw1HRLYbny
1nw/4POGiJIKLn8zMILlCHiHTnMttkQkTllkaMeGujtcmQ9vOuwc7k4IxEeeWyMB64VF6cHmnU1S
1yMgoanjSkwCm3EkUQ0DbMHgfhHY1AxmhfeeC4ivMpH7UdiH31BFh+SKwQbJZCx/nmRrDwHiXU87
K/al4RmQDrKsTM86RzeUSKZPgcYGRbxdBzaWrNz9ToPb2BODTBI0+wtQPWCulTYAW6xslSmBRsJL
0luNNuDOi5JVjt6phBKZ8o566I88iDu14JE7aXWq/6X7OcQg+VkXdhAVwsfLHPNNnfZm6U1U+Y38
ElG6stDM9Eiaimt/gvuxjtb+PrdIdQX8qulAwLM0G4xHRV/brDcAX9boSW+bYBJg/uKrt+3sPoGg
Uf1iMitl5n71WjQqTU5tl5EbRIjjbKarreeBP954X67rLFTr16jmsYa2axlBt6nS0d/Fmzi794VM
9s+0wt6yh9r+7IWbCwPnNIGy9vzUgIixkbfvc9IKuRiUr304cxre9iob4E5eLtsArMsIH6DqqzgY
6CqMKxJJ5zOJOTWUFxg8neO64L3YbrGK7cDbEghh1KRajapjfDtCV8ZDKXuPbeG35BTcVkl23ebx
yVPZ+yyqRuFWdjApmZi4zKvMXFIgb/lC71B+v8/EW906YZKOkj4HIazXSH9UR5U4W8/BdFap3PuR
ZtoyJUgRjZt3RKBfKZpcIxm6o4MVjvAadY85F7IuFZupOtg5XkRbnl34OcMA8JQzS33G1g1SBspn
u+Fdp1uwH9USpTvp7bsS55fRt1gtTrYmYRlaXxrRGrpHdj6Nlrc1Z4QC/aQIaTBRZX0U9owypwT8
yJtPjBNYNqlsQOKw6OpbTIdd93DKf8T40RJTODtf7JV/N4aeQ9nB6PCgvcmyWwegUm30jco/92PX
/GYoyBedVE3j5zJpUsCm4DYYnDx5GzT7CQCS7RhXwNLYRomCxv9UltmBX5o2QORJIFrUg6QSMsIT
IKUOzJJayTQ4cSnZfROKTfDvWyF/r3Ynz/byeQflOnPiSHZDusVVMPy/Y4IVCZx8QS+RlbYwtNDw
NYpjQ9jyO1bJRkVd46KjthYzi2NeQjRe8lpNSROYzHSPjzB5DXAYM33MIv+gsg8Qrxe1cpxZoZlq
Kg//9RbQemNYfpISsn9aF3IyYLmxnMcJ96TaM2CxgXKF94QXa15NOgofFF4AzbKacdfK7G1+d4Jw
4Bkrx2QUVfitiyLh0yWDXgsbOkhBa0j5M+F/3Wc7eL6Omgyu4SPMzcG0sQiy0CZsNICA+ihg2pwu
9YBys5qCBS6LOWHHoaPKHbNKooetmOhfgb52ueuWB9/pi4xmgifac9UGrzjg7imEtTvBOG1l7kMY
+csEwHwKtVIVZu+2+AyTpVFY5Ju94k4HbUsRvGkM4RYpy+MYCPm3z7r69B9Rz6JH87Gfo9vg1DmB
8X9qZjahVn5RLO+XLVK2XgddWOByHvfWX8PANUDzQXfbmcql0yIreUg4/6t7pIRuBrtpxMFTOT6w
kSDKOMerC4/MXdtsFqlyWH58+gVOO8murmhbz1YM2L+MnuRXwjRATJCyPUvmxzu8SEz7nbyvY15g
0c6JkekHGgcSdYmmrmuEfNx19jQ2Ih1h+umyRBk5LDurGm8GWM9M7+izZpVfwW4ElyA9AfEleVs8
o3AdsL3yxfTd/O8euO/csRDvLtT86NYO5aBueozsLDeo2Bg4WGoDyov7dLZNsHbLz8uaXvXXgpUy
rj2AyYzpHDD4Gmu4d2j+7MX7XvVI4wlsCK98EuNAcABK4ldJ3+pr4p+yFwI0cHuhZrejp9NSAk67
4FmTO1uz+pZ55BWlGl3vdZs74UGu/KJYEsj6ZZFFM8DGvLNpf714mBSeA0j5ry7BCizH5/yPtAcV
OKencMex2kLNVwn5pljjpgFtZsL2x6sb8G+W8phOpgflfFfh5P5T66mFNHak/Wa6yZN4qASx9iTm
NfNnJ4WtAS4EV0g3cxARtUnB3ELjJnIOLnHsWXB3uj3vx0W2SW3wl0nPhhcAPKhF1fQ6QUwUPmtr
eNRMiZzYKTIT4osbDdUzrthLRYt0ag/1MbFTLsrs2veDbLjY0QnUZCR5FcfR1RIoMAuceY0HN7q+
XP4LfJFle71H3+ty3QXt8wkvA17DnLLB4cmnw7nu7QdUmE9URyXtsiw/jmvQwsDoJ3Idzn0kAX16
iyBmyzaMb0wzReyXZvzX75nhZQJiqgtDkqD7DF611lkvg1CkIoIUuUyvncz0LFvZQ7wneGXVQPVQ
1Ozhu9OvZK9otgYUqN2ZYrXKAE35popYezoPmzFI9GtbXSIvcOamDvFVHGFN8bJHcMs2u4kdysxz
MKox//ZCZRIytaB7P7XLQttL26OQf2b3boZU1AGcuoNaqM8EAvJtaCpcWZbvbmRUiKT8HBh2CtbM
j9kvNsw2AQ0BMMBvXWMfQWb2ztP+KS+siOh/Ft4qZmpggIA/DeQUqbRwaWe58ABjI4ACdxhE6l3z
p1aI43UyHSEjmZ5bIzDoy3mvQZS19+4mCJzgbpw7XQnfc36nTYldwHQd1bd7PCAz3zTza0aVUYsI
l02cpoevq9WSy8FygUac60h/VfruKUbFm++9HdQXIWzHq0ghTcDKAZMYj89dmbDG3A78Y+JB6a/x
Yu+Do3ulhfA3Rn7Vq5akMIYOIcYpeD+GN17WS8ZVxNyKeWnftRXUZh8kHdhkYl4gzndIuBNdGIEb
IabBhwEI5ubkYTBluy3JKTX5jf7TSBIiQhgGYvj41BE08GITmyy9O5ysbN6iev6KDQOcDN8ChvIw
NaDE/pDu49EEavOGSkmr/t43VLolsTeo/+wljqfY23Jt5wLT3z+nyiaL3xDtAeXfxGhoK9+FbN9W
i4YcNUm1vpTPx1CE1mQ9ep80XwyFd0WATxutP78V6ghnoF1d0rhz2qddDTt0x159VA+1cswYXauz
OdLmkKsskEWRkc8iOpbPXZ19w53hpDNh2hWNlaWc7Cyd7+lJatkIYQjMUIQnkVkTQF4HeLSSSQc0
KVgYfMoBIAIdkVhvIMdUTgZSNj4FxJ6aIR3G6HvcEtSCtbL1Ztq5bW93jEKvrzK3C9FlOGv3jyaU
r6oDdLB/rGyg2NqSebPZDgo+W0qA7TSsIecAyJE+cOS30YaFLNmHU2+QzmQ224gtuav7EFrMWpcW
WCOys7qVI/MpqgKMCXLkpntvzp4ClQro/gQGnfHpkwjdUwaGFlLS85lliLdWk9iMloFZ3tuPNIdc
UCV3+Q5MoWHc7YcegJPqT355SnniKC6jOO1FqcAPwNJaDDfHhfplS4btiyiFeA79/+cGKv9RU+7j
ZhxCAEB/68nJqEhdw128/WyxodISsPFsykQsav4eXJ8t1aQNCz/shLM9L3FZPx2tBzQ1tqtO82ST
9GEhSAnM67ppaVzOyDpaMtJxYy62VbhDmy0wNQudxbvlGVfN//FQu1p2vn6PFAyT7VdBEibaPjoC
Wj2TotwnAC0IwYGyXh+TyeDbA4qfmD+QJKYo2VmbiQvBB3osq412DQo7Ha0RHbALOGi2InSzsLbl
mB3c7m8XUs0t6aSNYUix2s8+qJY4/pis+DU2fVwRNMeu0JTXVMTuo2qQYSkX9ZZe6DGLyBKURXf5
55VzrGMFKVd14aO4FXYP4MTItRPIVdJvOO9sPz4N/hoiso8aTb8RJCBGYyL6vwCjbmQkBpYIq93S
tdyYPaUT4l3zFI4piwi083dfnMQ2l1ZvJKYLab7xz/ITiYQYohmYZkJbD9kUXpx5h+RLwwuU7SmH
t6e05+cVIR7AjiMawGke7OMb4r6l1mX8n/l78KFLtH0HlNOlpog0q4U+aejqEpeO31QxDnGc2mog
tbK+Jyc/34UMK72F/SriRax+E1n9m9ZlykhrkGPebvAptf73Awzg2PNt2FHjOKGlBTQ1eTL6krww
18NZb6PVsS+3MKTy5V9EswY/d1KRFwr09r0cRCLMFaAV6G1dAhJl6hs+Ul3P+gsfb7fytfLBtaMz
4QRA+S3s0o4WIyIDiFLyF0NVg6zVcuC8WfgsyA1iqYoPv4803voCCih1LdoSBChr9+8QhxCqR69P
4tP3KubU7DzO219VzyiMfS5RmuJQa1daujolWTGlpC8hQ/7kSxSZeo8Fa/3uJEDxfTYV8QM/qVu8
AtRrMR3f9kWz4VsCSkQmHe84R9Qs85QuLVcrOm16vDo9vJROld5/vl+p+ESc1vUleSEgUnVg18MB
3b0s2CA0wrs2pp+wQ2Yh+qisN18/VMYQuQq2MM9CBPswv3N/oEXXDt5OFKL2nOsZuFwbWG0TCkcm
Mrj+DgXgIwF79FrDA8/8SSOwZTvEyJT32ecOBTwKQGbswTHYDo2947kMVeCMvQ4Q5wjl4Z3WZ1AD
LmD6agrlo4pjaCUHc4nwk+mOreDDnZ+ukDbsHVbleKXV8ys0U3CrlHKLmEwD4pRjueez1zDmiAgl
FoJB4QE3ZqoSFtfxS+wwFN+nqRQtpzaLaOf0Z3JhtRcmqTlLAq7dEw0zMGiG9UK1KuC8sPocmD9J
5FGkCM9TDFvLctGmT3GHYLbLzBrjlConxsLqxnH8qaueiTULD4gSzanUXIqY8G0zPCBaLmOu/97y
mkAauJkrW3nFsOCybET0h0jZ9/vUfQa8rlWQ+uVCg4N00KTwJwm4Kc3imSmdqXBDfgZ99I8BED/y
2Yexx/HfOGnMg9wNT4bdLV/P3xWxq0hQ8F+qA68zczzMRgpF3Rk0bvcUbI+Op6D8u5emJsklfRb+
JFigcIc578xxpviwizcaW0A4tRMcMqkENffnpgLV5z6pO87ImwFNWxkZb1/Jhtf2LPGGn73ozkTs
psPY/FF9Jm0dKMe4FUwLTJCf44a7kc5qGwjVWRrN1Liolaxq0EFs9DaiCqUYXiKGxTanhl7B8r22
acvvHfM+NFASL+44SY/n+Z/m33cDutelVN6F5shHeWHBLjq0c7KVA7m+rcbmA8pj4bUtpYAJRY+i
nK1+oOtmcdBJ0gbSx9XbL/78Bw2sACzj0a9r8fqlxQAJ4XFC3jZx+ywYAdD6krVh8MDxXEDBq7OQ
MvEuVdJj0pGT5IirqbQGpieUBXbzJybv0wGddQy9o5nRmmbSiuPTyTbIp2Uc8KxsPP37hKyTXLGm
us9xipe2hCrvnfHLLFwxuOYVHqxJSAxsIEY+rJ/n9JmZRw4SclLQZjP+M3n7UZMabqAjlWpRjykn
kSiTw3F+LFEtlT9hRoPuMmZ7/VaMqnOoE0rl82oWkGhb9qD52NJDMlc7Cg9MKfhUec1zNOCEHjof
bPfLHK7n+5x0v1vSOzClVlH7RiQzBz2I7RKiRMbfwb2f6kn4Aha6StuXSBdu0ocpACIQge5l8uGW
UQUEGSnmkF+8sDkc6UVSlukfOz8D28CCfOQptMDhtb1z/kAQgFaEC1uHZgAmoIb+LXfcgzXnGB8u
iKI5vZw3qvJ0VQCgoo0MGIQD010buijOXmk/trqqvlnIQ0sC2IeLDrkTaBPxIVXFg94h/jKtgl0J
b/bVM3f7rploy05gm50Wq3HwF6gQu/Ji45veq1kiOB3bovXeXikgxGjhxz4LFX4x1IXuezZf35Ut
p0uPI86lYb+HTe6iSvLgA1qoLxlo1uQzbWUYU4DFK5d08oTUtSHjC/CN4dF5W52D31ku2V/3OYy9
HVwitlIeXsLZso4XylBHi7aR1c4BEShtg8QDb97zZ1Kcg3uwRpUM91+x44nGzVtC+R381eYratQE
sH2DG82e38NRGXf1mAbPY6HDSAXmy+gLgNKUdKTEoN05BDX4yNHR2sFDuPSrrROCeolgs0+plfu8
pEPXN/R8a+E5KbBajYsYjHIEALfvgkdTe0+B9u0SD4cutbGmi+Y0Ui/qrLJ1nqehexxuGyUL40G+
zvcgIlL38hL7BIWrCyaEQlZMrNd0OCLmvqR2nO2Wro5G0HFgYJXYhX3n2vWVwLWx4HvkHe2NcRoz
31cUAOxQAllFHuJOmB2utMJ9RQbvG14tpQRDgAztL/KGyMWEQTBmn4caY2fimcombFi5pJcyKJYv
PLXO+6dMNuRz5XQGzghpSmXBbmuyQ60ylsj9lnzjqWBgcj9HfTaGvyxYQuCi6l7+ssquxKfhggFu
k/RuFPALyifGU6AV1ZEgEOLiCZDZwv57H8Clo9kcc37XAkgIEnYwlOwh47Pnbb/+Th2RkfVZOr98
ZP/l1hJCqpus0jleZebjubl6BdH/wZi/0Mm7t4QVHrUTcXr3HwjDDeb8eCP7d49QvmqVH5YQ4+6I
Xr1tt9DVNBoyusWS9x1Hbt+33Euq0dMA1HVa9fkqCLf4C6ogKTG5y8jOWGOkCSdoTLTErSCMNXbP
sIpThnYy1Kwx808Mg77CbXYoTuA0j6mlhNW3hjlCCw0dV8ViDAu+Zr6cDmY7dUtyKl4m+uJP4nny
O6GwOH08eJh1Dkg834uD1Dc9fDto8xfC7xpFkVrbpfYqackynwnFZOkRu5rHWCQqhrf3+b5W1WOh
Rjx/5uB9rFMTDsntO1p9ZC67jxSou+TryR12NWWh9npBqf+w6qEjT+DOvciepBDzqBCS9hAOprkX
CJeLp0MmbwOa2Br2CHAF2vSfbDvJQDNo1kzSb1iZ4BNqYqXGxSXR7SJ5WiNN/lrDpbnD7dFE2C/x
zPgZOtM6CFtULjU7O9liZNSN3CJleRnRjqnP78QW6z0DxZe1TCMC5n4pYb5gpDwC3XU9+p6THN4W
k0W3wXIHBo8mY6OhBTNpmMYfXQkWJquTaoTUGqC2AXLsUEjUNOj9Us6Eb6ubknaBN+vDPIYLEol4
HzUKPquPKQ7cd/Qx8xgDhB3rRPrH58w+YCV1zrgg53M/gP1y5+YsWSCMXRBhqxKHbV6ZAhP6f5xd
AoKWtkrgkLOh98DwH5Sp9uZRREyp+VWQ96UrHzY5nbqF5oYk/7JiULQoLFWbpbvSMwH7NiqVyTUx
JfEvVkyuaWXgkvpHoAv8SVqipigcbp1oFIIvqn8+5/9JdMNBova/k7OfeYrAusjsSAes7Z6RkfXS
YF1LWECfTW+n3weyqp6jhLRKxHX6ytqNi/0lKGbZUvDBuWdGllVjob25CsyF1La4CfHCzim5/fRo
Z0fHQKANQkStIZ3DdnXovNhJBfQ40LG3AWi2tgWGrNVuLAFZOJ43ka9r4WUNcz4ZRxOVCRibpmmH
JQpHCy4v/MfH9gSonSq3pVF2xlfttXJOIKBsZ3grJGgGbAC1qE/GtDl44Q3Q50Fd56wq+BQUr2Wi
CJxONqzD6dS2IrZvWcsY7m/RgiVBeYYmKYyIKc7eMYY2EOjlA0dKNwu+7GH9M6brmfAbc0KUha8S
iR9/djYoVzOk41pRWA80Gy1tQ0Lux1IpQBKlZyWXoGDnIQWyEKrX0T3MIeWKIUKmnSnfKRVHGd97
JSxAn/9/eJbSwfVaDMNcfRaxkQiyxQ6qOvrD+nFIOF70xwJOAZTT/rYEtHMc4w32npAvrNBcOqAz
7LkFCNFqlqovGaw+ApV9+bBaRKp1bi14GstCcVIdmqo0O1ngHWEPH2wIeidrhrCxJKCygGJa/cfq
iuGAgpoMw5gMU2UzoZhKs2u0KvJjpaadBaed/BBXVCKLk3ldmLfrcXjkB0MFa7xD8QyJSm9eozhA
iSahOsVgHWLUxG9b6Nvca+8XIiLexqeb5rvP+N3NC3IXvprXWGLYiOP7o2HnaKkCKnZMao0ZU3ko
Xfsk9IqTiCspko2KrVPbgH3pO/rCelpATBy5f0qyvbIVWJCrUNI90r6kHjsdjFKkgnKbjoIq8Hgs
C2Xle2qsQICjgQzn2ZJ9NYDv+buZyGnDhxWjGcQ16BhUKfO3xa+iBHwv2gWfPY+gy3Fv2WL0TqNx
AWa6d/UOf9y4LvMTghe9pglRYmj2aQ37LB4BBve6ftwTlWu0U4N5rrAHevAXwKGXowiplErayABV
7zdC3w7yoNouHimQLyy6YXMPGPmIvv9aXGfff62glV6FUOFdbXBK0bgthnZjN6yPBY2uKNUYS0mv
ELmQy5fyNSFtAZAbARApeTqP+ngW4L4Lw1C0C4qOxTI0s0JRMD/W7wk29Vav45k3m/ebary3e7qV
vBdxe6Tgt7O24bBs2krHxIElfYFgm2k469K3caYjL2M5mZHeeJbEqjVp/34ZJl8vRD3yN4f+Gwac
2VwPJEgg/42lN1KUSa0BY4oznN07vyi+AfYKh1SWbb+w+3QK6aHqrlVgPCudO+Cj/HgGyjNtDGmM
1S0cZvGZ9iGV2VU7sCazgU4lHGcbP5WDPytndLAWRSraALv2/uBmdDm37GgDy9URfrEQFYMpRDPB
j4LaO3us1tp7pKNk1pZCzArLMH92RK1NkxGhcFQtvFa4zqp/jl+ajoRrPmpLvVJYlO3+qTAkzHF6
cOY4DXk+EqRsleLeobqcxsjA072lr3U87YXocXCpslmVc0hk9/9dC3/OpbntD6Q+0lnuHMKSxcEP
Zuv0gYpkZ/jJMit5Ci7alc4ju5FOrBAkzkYv5HJqbzvv61U+K93bXuSyIuNH7pJe5isYN1JaYq24
wjp8Lx9F7HimxtR89DF51rHc1Hm1gVYcgrGmgONQDqwwljKJQg7HmnG+OwwHpItY0ndhV6o8+Fob
ksHknHTPTGM3vdOoiNPKTaJJS34g4jAffVl/bbzR+EWNaa7n3+ibHUS2N7oN9q/MLX7sMHrkuURv
2wOdDz8zrga1DulQfgrBlsGYKOxKUINdMUhUXcPIUqv6/cdt31zp9t2ywWyfqD36V8XouF9Ob0Aj
cEZYxaO2IL0XcTUcecAXhUjivgI6JTz2E1mP/JRiFCQPRKgd3zdD7DcFtQ3gMniksorcBhJevc9H
R+4D61OAQvpLjwChVgdoqQjyNIcLESXBBQiETxzNo+xcdIx7oXK7v9VqgL4z44ipLJHlBTutOm9r
t31oBg4gh+VoXIFsfIHlKAWppNt7fBvant1iEDE6VP9taRRLUiN8fFJ5K40XFGSr4gyTO+kBf7T6
naLpP7aEOpekOs71SF8cIxV7kheDDsjT5/MgyRoAFmjzWWaBVE46t2+SnVrvvtczoNZ34jWRUOQa
QW7rkT2e0M4bFEsz+h5GEn6qoPTgEstr0T1CMyePo/bp4d+/jae0Gr9Lhy0CTQFmg4EBkzBb0Byo
ErkzFB43GDj5mf/+6SNiv2lW35lddu93hDIeo7hLXA9WhBHzTJExdl7obQH/vBSYWYsDKwRsR39+
0u6zNl7nL3PriBDc8d7gngD/k3YGVm9Zg+YC5tFwXbu5nE7Rutz8gLebk0ttVZqcWXs/YMfiOiX9
5pylyyt543GGJv60Blu3+G4+P4Lemo6J5qhs2bGUnIG5fFiEf6vh9A3NslVADsRqtGk9gS63lC9H
qEEWrCcbEc46gdAgNoV0He9a6cNeahrmqyscDSMbKEdD4sTFcWw5OcjXKN8MhR7vbdWG26DgWkJZ
yVRL1dCVQV60iNP9i1gXNZp8jrdCcA3l832OzN2VbhsmpC6b2xEgVAkzw3srXwkwO738LM/GcqKu
0cQcwWPEUdYlcFl+zzVeXNCcLdMof+Vb1vNMKyUeIbvP4P81zDNu/0ZPNyNeJNflAV02GrTMon2q
iuEyzvOrzb9H6YS2FmyOr4nC1ZVDbbboIYFD087UUGNntPyBK/j0fuipCz1W6kQyxP2aPqey1Pbl
WEkcz7zGviNsQD9157XQjNj7k17dSe6h4DBmhJ3L+8OpWB+rNnOTZGbULkbUpdyt/CXh09gjTeIf
Brql60pqm9oE3qXlMEOYsZS5tkURIzhLemkMQjOQP5RXQRiPleGmpHyQHRAalBcmlnBeEMq/PKGO
WU151uK3xmgrpx/GhrnDd5x+Ff5U1qQwHDKf/p6CBYuau2wKFatj82v7KDhRbUn456g4j4/p40ph
XE3dkH0GTYababEE+ViycGU0mUpS6LKNFvcTuiPfE6U2mNZQzjkq+KRy3vj+XqEmXrl7jDQUq6r4
d/4yIRpgKi3rWvrWD8at4UiLj27sK5kron2W6EECl4/v/5P9Rji/piRoZnIgOde/onBMux3do6D5
OATD8vI3oS5WuUK6CutlW3q0IZZI1oh+2RepAwvncyhRuJogAhqeA8RvAU2gd1WlzC+usY5M2Kn3
pzWfu3OtyPkWwQdgXeOtxyZLAaB1LkzSTSZ1UP+9NSI94cARSsoejcG87qgD9J4WEtShrwPVDljB
J/rcwTTJoK9psa+UN5bA8wVCrZwKFg0swa7e58qI6I3cCSdUg3jog17ct1lLR9cfN4hLelRdaUhN
pGW5NGa4mxmYmtYqyfWRUFEUBWyFiAhOpU6IIpzNBBBgC3P1lhfmD9Khhjf6zmvrdyYdoMnxt/po
8qxj9jh05RrPxT5qvo8Po6XjAczWXVDd632/hgnoVSVh+OInjTlNuqLf/oWtiBMLSWKe03n7vOvK
Ae0zSuakRNYoYH1lDGNpd1nWC8EyftvZC7awVOHNQ6YzW2KLndH5+zjkHo1J/BLDWBRBRMdaniZo
wnHSEaAxy7VYyoljIVeHDwQ7szG6YAYNFKaH3vjuOM/eqAP+njIHgikmAE+zLJX3O0Y2d5sduZX4
g67/yVZj/Cxsui+Iy0Ct+wOtdPd06Q0W0FvaQVDY0K89Jw08Y/HFHRD/yl1p61a/qkUkMc0i2sfX
O9zj6s0MCuRFyeuJ66+ybFJDtwh6qGcIK5A+FDWM8w0vi2h7H3g1ymU0g0Pmcuyj+LkzgcahSw2b
2kO2hhALJWWTBPz0TPzz51Ws155BXZdS7uREebs4/XV0A6L4PkQmSB3M3y7sF9aU6c0GFcbVEMRG
7KzFRKqNPofYAb5PfY2+/fxCJW+T6Oj0xq/MmaktQd5DJwMSAzPnzXGQ5A1Y7h4rl31VCijWCNbF
gsuc0vkogRvJgouNcKhpXsjA7NtlxozZoEGX89ePIKnIiS/Jch3YZ96tF7PVDlnUGtw0j5YufUVy
O0uwnst8pw9Xv8oA4sdOqJu510ezhL0MqiL5kcCJEZyt5LrARUjbKmvvrXFbKTAmft+HdKomYMwP
OR+fTaF7IuXw/60VGXBYChdbwABKqpJnXli6jk00GU1tTtOHjVypAgPqjfxRAfENUzHEiHMz94VX
6wt3g7EOApm7Zid7lyCCsU5+tPikZVHj29B9d4jNBeW4qTYI5dnQk8AY0+sWBNpsjXSiwK151hNv
J7s3MeCps7+dErsrKf7imQ8R8lPNsiNqEs/Y99rkz+SFZzJ/pEHmfEHjvkioDHrYwQ0E1Xf/rywc
wf6FdXdYdT9V8IR5JEcCzEsoVTMxVAOJFEmrRPmzQE7ELHZglW2ZeVqUmtQrXblqkUrQYsCoe0QX
XlNc/+3Qw6gV+Y9/aeZZGAXCFfUN11Q7EWNEvwGtR892/VDx0DFW0ZXvHifv7xDaznu2vW6q72m/
afRo1+dCwxRVVGFv041qmzCZ5U/saggDRunhwpD1+pIN2EqvbOeh2amg2aEqw2St4QJwBZPcdBOS
GQI2GkAqxJHDEuHgLu9oi8VTV4HciZRENZq3Qw5J9IfphPOHzMcESVU+tf7LjTI9o7cyF86Ak/eJ
SwyygiACxvOLOZU3v+TIqeiY0DOMupk/jgECkFfk9s0w8/5QvYZ5kLXBv2kscIspvO3YqYI1y15s
Qgj8vaun/lOAUHj95xpTotHd5/H9WjwK9wdKaE2AzKiS0xBW2tPiPLtM2BkmdTgUOK7+aQZe/NLA
wbB3Cr9rm1sfevYGMWZq9/I5bNOTFtoMuYP2m2BOVjV00Rq9kilm1+DhoLthiaelaxIpBvKEalm8
8xYm+dPsxPYY2x2S5f9bKVMFiSGhVOFvg9KdxQoAXsk4CSNp3ReRyk9LDVTqth+FT67yAMlizhJV
xPA+KI7BGbnDwoT2XnTmupYJSlZCkcybterLU5tk+Y6ke2Jf2rstAUPG8gLx49AgNYqP7wKBzcWJ
I8IwsXSrQntMaeeqzzk6nye29+ayLjilAITsm1UrWuQeqDhFevGr6/5hlCd+EQfCY8kGL8Ld9Of1
j0nWoqjW+xRcG9H8m0LmIfRHpDA7M260nbqK6poQ81BLmASJPNfLsgM930ixcDKAMeWnjULj7sR4
R+yNDeTr7kxwbnrUVpcbRZS5H8wgV4UvEeuYtc6hMt5S1cIP0ubtvWLAaSOAGD2VZk9KB17hvpRE
5x3p3tuAVaoZZblDU85VMXUrWktegDbOeAfmY+OK8W4NGyHIJ2Yy15FSi5YqSc8cisF6kOCoK6ey
Ztp9TW/gDfqMdNa3BE9+NQ4peyphPN9kZgUts18o/VSrawu70TgvW9rfjmHIaA6QjztPGfL/EXcy
4ZqVLHKpdgiEuGKeT8cVEawo7O8iL373ORzMZEEKTbmIFjob5YRughRr8IPAFIgQdv0gO+vG/nhO
tiNEl3Ds4D+SabGL+FWgIHuXJ63+KRZvTD36gi/0V878oZ8BPF3YcIllFOW/ZLV6BcXW4fZT9og6
n6D+PCr0H2VU4epYfnp5eq+G1jehjXSTLl5Qcg0AvvB+co1NkLyB4kJ3UaSp41DfIJsR4l7eqA+K
m/HJQV6VqgVI+PZdC3oPamEETQs2A5pfoCQKBlGXBl1NIMoidmiACUd8ChoV027ZwyGXFFRYFMzE
os2yVjX0OIp+aXS3NI4eDJvBERsJuPTxbse1p2P6nrBxhr3CzuW7gBtG4NsCmH8FElnzII338LSq
jzp0Q3OUf3uPfBl+V1mPMn0xM/48twH2EEdzJ/eoovF+DP5V9NO6QpK0lv26JAJvQuZgkgbbJP1e
WDbi7F+lSvNzUH4jeBr4Vyk2qDenU83KpeFbBuVPBH94zssYjlwZqeRFp+TXjPuV3KE05Sws9N45
B3xBSgvTzzJI8Nmx6ZtEDLCs45PSEYny/OKy8XONnGszF8irdD6Ddhkd6HMpHjRKMyk4HmFOvrGg
yvE5bgfQUN3+43NzoRb/QyOj5zOjFAKSTNAeexQRXtBjHBC3QaL8BShXdj7o/seWG2pd4UPD6yzS
dX6dB6OEy8V1hSst2G4zbIkTzizdR+UNkoUQXMW0jgJ6K0LNhbqksa/wVRvxM08W4Ub0Y7F+Itv2
ynooaeFli7kTUyxuxxvDpXwcFGb0Spe44onC3aI6/VsMeFkXwQI2vC58dWk73ZqJGX4uKbHwInkX
Rkpdm0tRCOUl9GRmPb5NKfraS4e746/Gal7TRNivWupj37EesujHBIGwbhn8hOtI88KlPi0V15yE
SgEY4H0gCsJ+H15ADH3aesseplLJI/Eucyk1CwV6Z43RasYHpJOSO56YZrdjTtLifbFh3nE+pxPr
EJrYOWi7MpUlQnOdUW/L3VUR5SeMDY++tn30HlRbkxP2YbM8z8/UvTvB1ZqM0hUDsByvRXZl4wav
+1xbY9xzQmmJBtTVFLyTRQCAkW6Rc073bTeZ6cs/1+tUDE7nN1+n1oPp1K3uqJEV2sQs4zS6F+bD
mo5VafZzxS/Ey09otuXW31Oud6J6d2MK1h23QlkNiLae8w36438fxvy465gtjNEgeNkjr0j1esCW
perSo27wWoJ09z86JilugJJLIDngwA0KI9X5UTt2xw2d5J3bpXj1lmdToVuRHT5aKua5YM9FS/6F
kGenYsYYLHgnSk0jL0a1RuUK0L/Xuz5vTe+20LXSK1iAy7xz/xWc8hjLH8Sd3DOt70i4Wd+jWIOb
8W/q3WJ5Lubo+Gq41jkosnGNIxkRyncNfc1J99QGomz6VpCzPTLvl1HoSlyrOiw+ef77cYgDwhpt
KT1DvRf88a0Qin5CVXX/ZvsiW1DPbZI6GDk7sVb89bTNo0jvtqmDduw36lFGHnEurfVInffKyHsN
ySKOO5GQiYoaImCSvrCvas7i7hIHst4cKqUlWnG2i8EW6IhIdLcqi+hwuPtPOm8kt1OZxp1wZuhK
kGzTvzI1j9JAKQBYa7dantAPZB2H3ehrUP31lsJTW+eTk52o3WUfJ7GiexUun9454iBhZ9YDFIUA
XxtXTIYZB+Zu8xF9xQhz2KWbEIymDWZPvsYF6oy+lON6YaXT91Xvdi1nXadSVRTtUtoubwiWgYwf
Ejt3KS2pyZIGJ7Dhbxg3RIQp8+uO/0IqHiEOnNmJmTS9nbek0tFlgHauRh5BzRtztAc6xxIt+UvQ
xyb25vf4MVtiAbL4xaAkRNORrPbQbUt4CL8FKIb2+b/YXWOWBh26qgkc5grPafyYZhFgXhdm5aJy
4z/cxn8YODqPi8Nn7AuUpRv0iYoych14W80vwIMQLKYpg5lrQoJ+7w36hEoeH1ka5v6isq4oMsdG
M3Um+/YXirsyJ0wZcC0fct2vYRYaGNKZeMAWKQ+NXtF0V5o75U/OBZf7BGyM1HJf0Jkhck4rtoVP
CCR3b6g9iu19MvhU4zlSgrPcq27AzeQ0vfXKn5kM8LjJju7moXg5nkYTaV8sELhYlyT6x3Ib1wWL
rSLOzWLF6u6UMYnbpJtvjomcbV6EKn91M0qRSbPTI4aLNJts8+r9lvNOibRN1miVawOKwLpGlV7x
hWmfbu9p7kyRdiPt30B3ECj+jlf7JW7hNBGwMj4vsfez6CGr2D3CrMZL0xiBZWdKHkaDc5rgv36i
DwqbrB+h0yGq8nvY7B1v8x8WTBRUu41AAjMdYpPBmrUHIIje1mb2NvaS7scJJVryP67hCPl7aSIh
Vf/1L9qGQ3ErqN6X5Z4ii/YP41Qj84G/8uuH/BybEjE9eAGCP2Gxx6r4XQKtx6tlQJDCto4DTY+n
eJc/5liOwO3icmEXAp9kGfofifUqtJeujmdc1FxqExKvKWeQPJfSjg/aDH7Hux1SfqxkuE56Ocsv
G/ajjdizZn2Ki9wWUCL3zc7D7+iHF8qyF6Stq4390+T/iASrEdpbiG6NzlEx6ztSPbz5TQ8Ku0Hn
AoiTeA6qXk8lfvkt9ZoZ6QifKDbDjUIGUtV8hcfsnKFwtEK0RfbF/+vtKaPmPlFpEb4WGrAohZo8
B0j420q+3zxW6FFmxt5N/2HM0RbQWEk7QcWqyqv20xf5VAFoqh/6JCzSNPZgZoipCNi4vf++gqR0
9Xd70XWIKwuZ564Wg3nwmQ3w5+EJlVfIkjb2nOTV8r0IApGSiYGvKzfxvjDV4CYqazhoM2VNGxr5
eB9RIZNVBh7ch8g80/T6Om/ohoGIVI2RRns8oTNsJfWSWIsHOJw6PyirbOGyc2Chy7k8EGeFMvsa
msHrhnrPXL9A9UEYVJ9A1XofIOS9192n13qhFP6pgQGSyNMXBJyvcOuIubOC+02W43/UAPGbDAbg
mzZzuVu6F2W341jSouLz9cDem/dVORRQH1s2A8c9atsK5AkHbUtZrQJZTCUi94dMUpxbaLCUvV8N
N6ceOfFoPvvp3XfKMHQI9vgkPSdz4xHoRef1Bs46GF+voiPhtOBAqrstt3JnHveg6JOM5e66ll2I
L0Zwn0wDZAtvOSoCsdOxyfYJUDBdJ/JTNNssvUn4i4vVbSxDo5CCB32F7YW9Lkf64bqXOV3x0R4Y
W/XjnzWKKCwWSsrHxt9Ej3XSj9954WcqGX7E/m/pI8aSFLqeKt/gh4En7U+YdvBtrcjTvwTtL7+a
3606RaIpW323zMNdrp+Y1t9NDBHCY5JtzBJzzeeXDaeTRWd6/B/WHG6uzuZfsmq3rbOx4srr3b43
7jOMI+y9PxSSBbwLUyY5m1Fb/AESKB9CdSdh4D5onC00ElvM9W0Mgd2gJLMXCohoShAWbLfu9tYi
xsuq1Orm7E5Qtc4evH1aDQ9a3IDCBH/r3da0mq/YpKBAqR/d2yyoZaQ+zwGX5zX5G+hAbg2HVFH7
K8weFw0NHf/1E8+P3yAxFdoxVo1U/fe05v4za+GL48093NploLqfAqDmyXl3VvfRexwlysWg3s8g
CIGCWq+ynooSth5OS6kIKt58qtdrdAPsaL07zoIVn0dBx75ewcJIDap3znWWCGx/6olLlE0u1UHR
fhKnp97xvYtWZVZti8905SgmO0Wo7KRlihSR73AFkbz8JtuH/TthALwWq6rvYyEGiOTSTSbALhnQ
FwRWdPo7LPob6RMb897EBSnt8WQRfc0ZFVSuC3DYnLpLO3xTxgpj78P5UkJ1tqfeq5nKy1lfbk+s
Nk+CZDNJqaC80coWnomwozCZwXthzA/48OlD9lmbtOWwe3dOzIbpKCroJg21GoxlsOEq8rn4Elnb
jo9VRbv1v41x9JgLG5XjhhdtrjA8JRAkjIJ1AmNIXA4wG9e8dypyLzkfdfy+sWtktmAV8DJELAjx
NYY4GwdILJl6I3dgBgbgsdO1tQMFIrenerl+ubzlCior8ahpi21IBmaPwR6V0MFmRs9miUEb1Oin
n4oCctMXxYATrS2G6bnIPIfKxqInm99uoZc4sf286o2rx5QglXW5b5AbgkTl52GfMxlNnsOiKz8Z
nkwClAC0B8P1fBMOTFGoSCP3BfuPKcAHSHwOHuwzV8v8i05xi89Z2xY2qUAQF9kGBZAYQocraGIG
U4eQ4DPwvYYB/KeSusYpRavMLAnHG8ldo9Me81gv/UcmsssfatJ+tidIUdzcJ9XukujLYXcs85Mo
obrnVcltoBm8I162ezVrqCfHrT+33vMJfIsjdIY0cnbYJe80DyLRKMAtqiSVwaq2oww8r80Omshe
1CUU9GpF2qd31yXtJebeUnadMs+bZ8cYemeQoOwuHdjwEJ8BFAysYf+nPwJ6vz2DES4+TCKCkTRA
nuEGOsnscijM8R+Aug5ALjWQtf8WVy/wkN0Qk8G8K+uI9Ejt3f26zSeq1IZEkOb6h0S3IJ4VZMFY
wUg+CCR7aAgeWWPegJl6EVkImKavD4/WYuDI53WE7sRK4FVTTa/szlJfd9+G4J85C+jpccO2QZ+9
ghCZA/0OL+vZhVptf5rYdxwyaD2VLZUIJ6sXMwYxrf2AvvedVvXiDbEu+XlgtTjLa9v541bA1l3C
apJhk6f1ry8gEyseuKUDJndxkUQKsOvbjyMqq7R/RJwfwN2lIRPHba79TrXQxktA4aoMZ1HB2Gid
70kd3cmm/WH9m70xaDhUqjRjQf/cfslt8+jV984ugo1CRFiZgz8u3mNWSiINvj+cSKWvHr8o28oN
j2hABEM4NvjOUSV/M50xhywnQe/6GM7enc0alJIYkSzAQfqM40jW10iGwdNSnc8KXjcT89x1Qmjr
3fnR7KnGEPCV3QIJdVmIBzmYz6BXneP9Q8yfVTQ6cdJgu+PAhykD5Y5EEXq5Gw0A8u1xbXHROQTP
wa1icItvLnDNQXTvUsuky2tNJt+I8Uf3rVtZvp1pAy/H9KhZuC0SSnplpRVE2d4gv6BKohT0KeEw
6ylvvrlvknotQprDO2v4e9jmj5wO2MTl1Vd+P+K1kRuQLKW+Bq0dZmFx9Wm6vhzePYAi1iGSyiuN
RQfBnsnOcm5bQ70okJ4RPhz9WZOSzOG47INoK4Nt/YJbZzuDc4tWmUaRj3Fna67uhkfEbVHaGDiO
E8KXrPrkhNGpP0bCDCEk7YkJC6vkjUyPJ+U/UMbYkudP3K+VmYOxID9G9yFMhaRDB6tIXvY+cjsH
R1DzoEQopY+mq8DiRjTBLJW0vYvOBLseFKBXgGhfM2LFeh0fQHDYKmkuRgmyQ6Y5vR30AWKtRFcW
r1MChqsUsEnTAzswZwvF4EK/tq58fz1EL7xQDagA84AkUU2arzCalbeUBQGFgy/DxCRQDFDOXrJX
2Ampa+Mawevu2aNgYktBr/UA+YNfTexl/KKR6sN4vCh0tvAKmonAQJ3zlzql9wYXT57WpRTDHhWi
ZrJMuqm+NKY7r3BmxkDFvasuAXEtUeEHf4AMwJrT2Imn3lxQ6B0rO4T+ZoP2TjHI4f/nxPxsuXeu
30Y88JoA2KLBkJZ3HBRczwbU+X3cefcSa9OZtY7cEV+xbU8zmQGV07NvC82Osa5YU0KwqSRqOjH3
Kd4f7U6qnliqFXiTgRq2aovHPBsPkczMshA+/CqypoRm30UZ7oNywzF77Kt/t6zEnU5oQI97Ymtp
IRshtwU9LNGS4FlCucsFsiqr+V2OSTiMHnMz5WqmVAk+4oW52sXYK4bSG46tgrewsxspOpyErm3T
QENqHyKsYfS16inpPD0YJS2+hjudp/Qzepjf5yaz4TI4ZHdW4zrk/GKrilXb/ClWYokwEf/LjEiw
VurgjdiRoAlJNB/VTczocQ0C0nbK3FvbhATvm8JkhJWONsRa4UoHk5nBBTNdlBE0ryMZv2wUdBEb
jZIVNVeGDtyJpRiV7oKP3JCqGUqm+ikCSv6TbHXR1fK//PvIPlUqChJBTaA09cuyoGbjfK/XyJNk
OZLwTc9Alh421W76vsqBh54Otr6GAUPiQ3Pa5Y51ZdU3kuTUrkieZ4gkhyni+Cz5zg4j9S3Bb6ji
by7ZiwH8U5CksGpsX9h3JSHytm1R06aySSTOv53oJ5PCJWXnB1aMiOBt/ptgH77SBsa6I9a6+YP7
La77QIl4VMdORAZmHQBShcSlOkugjjayTcfktuiq+WfbGJEgC+m/U5dW8jjHB5mcVlpcvwWnufvh
7WC1JWkhyvkwdin4mi+HrlpTnIpI5Cc8bM3b4X8FT5RNgyi41mYcY9FXBOnSzdsjDaK+ldIr88zS
NT6bct7OudxGlJU/uCCRCSplI1MBPBDbmOITUWAkGR94ComPVji5d6gfAA20sgwa1d4Nj+cLGdd1
1qCfICv/t3koiOj4KMAvfxaBvDeytohEYXoBce9R6or1oo8Wu+6gbT0Uyy0OxB1XSz6MYzip1R06
JmqVSy/EGww6wW1my3yjZiYUUUQkNe1g7pWq2jveocZMxookRBwwsa8nGqZ4xC4gGPC14b9e49WO
IG7GLhqDTnte9lDZZv3XyBu9UE5Fw0+FoWP/whsOexjTkSmxwjIhXw9PtUr+KmWtu1uCcrtBp6yg
/P15Cy3CvTzTm5Fsr0oMekiP8Ql73ZAhnTTENMt7FywzEiLt7rtHX9cLErGzwdOJ11Rsfoxb5ibN
bTpJ+OoV9G1ElB6RFuEYLP8PIM9hTryAu1KxpUq5I1h5lC3ncUUEUusYoQeB84yNZrpX+cZQCwED
hANUWdEkPteFCJe7xcypib4k9GvlXtZz0ZzLggIb2Ob5co9T+xi8NdVxbM6Ne2e/fEDAk0AVHuXz
Iml7dqVNvjZXFyjJSyJ8PXhvByCMWTosABzJSNCUHD0qHH1S4fHSA8em3s1eFggcC0dUo9v4hjCS
DTCx09Libld2E4LpMLxHnZDliWHK8ddTf2khVkY9BK9TnGamWThTeX7G2XDL+bcRtKT4nh/JCAgc
tQExjQJp3siJFGcKnTPJ3Qz9STynzdatGd4MMjl41RfaQgtrBGb391Zt0wYFS/kaJCAfCqJ8cUzF
YYrFNl8allbVQfQgsRq4g1vP01Pd3yJhF4i73QvZpxp+FfOOKOKxbdfvNrbeKR767gJTUBmleaEX
H2u6kwe7HTu78lSj3oLlB/pM6nqPzmsYxOjpef8GjENB1tW2Q73zV1JGEafo/a5iP++DgkPh1g+p
XALdZR7j7HYRR0bItWfux2hVarony6yqtCdHgXK7BhzzzwuX2PfGeQIaeEtB69JhlB/5Av/KMVCg
eXpQ0MQ7VMhXh95qlGutXqAxsSTgmyrWagENnInmCC7ShmlhZ0qGnP4mZ0nw/dIEc1hMkEIgXP4X
yLQIqYYhn3dV9Jp3/qzmQIVz2/k8IpbFuZeXMcq1tMHIAk2rza5MePs2BnRG0NfRFEk43C4BujZl
y0KyR6p72OZpnZ/SbcGE6cy0dIwa4iA9Z8ODS0tGo+pCkUbkKuXwXnocifcJ78yBi/MdZLvcQaUT
NCrLhJJ0gTsNJyjj8SR8RLsQfMXXetHIKd7xcSOjXTo5IW/uEHDp4y6BzqnUEX1+eE2KF3Z+V9XR
SPK6T/KqhVFd6Gqot4dxsaBu+vxf7Mklhd+NbWR/HgLtXfr5KF5ZpVinIWd+vBcSB0A1zkBprOFk
hLQSpHRtrd+mdwNWRXdTU74pIew/7mitcmY1joEUFhwU7mu78Q5FX6Dh5rYHp2J+ApGKknW3L5/6
FEcuv62IfiWut5nr6s4vEmSgB7mxwTB0le2Y7Z+zrqXjTQSLeqaBmsdAE+zpTki6uA9WsMks/Lt7
bv5ZZXP5XK/V4QEUbFiNmWnfDxaIa+wZ3L9IWhSW8IbPWurDxMx8SRM8kyOH5uq4J1LI79WME9ot
BzYkF91B/95OgIdWfI5OA4FwtGuMUP7aZJh5lHgh58ZlkKO5L0JlhQ4w+QdrQiAFX140V+bORMj9
uUB2nW4Mod4bL9o1XuGOtJzNGA7NpjWBiXQaFfxjvlL9l2SdrIyj6CcToJPcnLtkwBvOalR751us
jhkLSjQfONOJZLNOPRrXFEMJ8hrAYBRp++rW6mGQXuC0S1vJ3+BEZMVhgRK6KX1wZ7YAoAPtK7Ud
gRK+p5s6/yjcRPTVUYJaBh5VYnPFjW4t2z6IWQSsSzdkrEHvoZsV2l5EautTOW2GNNx2vYMe0v76
GUjSYJ2tiQYCYJfSbBmvjewSPjIjwVqsbCwOpel64mscXiJJXV2xPjeZbKIa7aBoIFU0d/3YGJkI
+3kYrZvDY/tYLy3P57/Juf01FP6/SYFrTeHcEX+35p2LMis5hXcIkjsIlITePmy1Fga8kX6qKsXL
tKPEjZMS/xADCABLJrerif6MEwt+2IIFh5AT3KBmfDwdRX1D2RD4w2KL1hS4oAg3huAbHUy65gKP
7tG6d1ev0QGbDIpcHXIRzsGTeE5In+8bJtMK/Moc0iPfWUtI5LQCh1vuZYR2a1Oc0wgMfrf0QoSZ
TfbTEUwSSTyvWsmj5gFDSVvRCUenG2zfjOj9pwFmG6LTWaYNtqUNKZt1S+fVZCMJcTpV2IAifFto
4l96RdYWAKdyfkioNyHMAUK8f0zszsZ7/QM9KoToRs4kJnN5F/TJ24+EKh2BufadqacZ/t8HSNRl
Hgn3gWTIpSmdmO/zc8LHg0kWWmKyLeUqEJXZ2Xd3rPEaDSqyDubeFveXQOs+7I2O1vV08JcNsZzS
y64Fz5lvD/yWByDB+jiT8MG9vRahp3nAqhwgC52oWp/7gTuINTURLUM1EZEdVQunFQAA5CM69GXI
hJsYMdEWC4CSslX2Zie2slx7HQMi5T1Tjns32xQIn0n5kNXQyeUV0K3HbnlHjblHm0LIDCBfh+lj
uU3vU8G2s0cU/P2Ix0MkzSxgE9T4pN6VRqHzs3kZW3MIk5hEvJpLBGTus/AoYwYy2PAXFu4b4UwJ
X396Bd1wwfqteV1JgxlL2OG9D6i2jkhuDban2UjwW6JhcE4Z7BzZNVWZtfJfltBfVWGw0BqGQpCs
tnEGYBNACsIqbSNBK8ujCMPrKJuI9gDorFBfvFqHgSwyqIOt/X1mAzWDj9oeatdstm+CLNQpbLqX
isQo7uwH+QoaGeba/aizTJIXOL5WPUOJAjA3dnW0Kqjq91I1yspUN/xfmDYwYaE/Zkl8GkuUaGE4
/X1H00S9cx5Fm1Aj6maa0NbmxmRk46UbEbUroHIafbYgbw/gerMyNv+xPW51WDOTEYB76/ckHICi
so3Iqj9UsGRullu0rmbMa7bQ1xskVSSrgovOLwf3riNcdqzatLBQ6z8VMG16umPtMAE/zdirw1QM
6EP9ROcAUxGD42mfusVuQHz7jgJVXa95seNiW4Lh8ByEjoIRtbWbdX7n9Vf5TMAxhAzh/l7U6Y0k
u/G0w7EUvWfmz+7Tp9ohLvCpp5SXFLgrLnP+GGWIGFRWnus39Rog2rY5Mc3XgoD/vMJSKIeBzH1V
AHP2ZKfVxKbfvGzkzQO5XgmEGHJvJ5L804LrdUHCBvWvmOgmdbBxH7JjdH6XtF06rRp51pQXO5DL
JFyKbOfEyPScMjBcx4WXDtpEbOZUpZtfL/BN1PrNDE4p/C4kXMTPB2HBg9Y3WkBRt7afJ3Vnxzak
zNsttjzY5Vh6VvGaHMc2eRrjJ0qeffwTTQOmcJ3olDg8VjABA93BJq+rPB/4PrY1CI7F1nRLCC8W
JF8iqYv5AiRyXW/uft+08P0ux6vuigdkarpXa/Ip0tddHHq0mNUXQW4Qc0i07H2+noMXWP17dlki
CQ6yO2Hx2gLKRBnODQddWijK39BZCnEMnxDjvlgyisvr93zt16a/ayrlonIdSBiwZrtxZwefyb7g
vTxtH0bh/vG/dcFh/oc8wAqzo8McmNgK7vYJk+rIInh41eL0zUUn7p1s9FI6m+sqrb1hXDLxlcLj
9XoAYnZbw1CGzmpqwsVZ9Ed5mW6Sd49GwUqNsQeuzQu3rx/XCFzaRJlBxYHsblkBdyrf9RPSBedw
TOjCdjSz3uGebyZwsXyG8OQxW1iG54Dwf/BQ5c7Y+ukutGEAhkZ30md5/kDgANc66iZyKlDy01eE
XNOokgwyQWURZ9Qzb+eDleg9IsayFJn0rxxTVDLapC9x9f9tIj5OcnPJ+4fsTBmmcdmnCpRccHZ7
f/zPEfTO2b2AYDGx9QkHgIu3kGoQdXJV90FesQGtd7g7dPmMr5cmkQ5ZDim7J8CjKG/xg8b8lV7n
ZGJrc0rGKmAh5cXNIiFkeMVc+VkARJoCO39OsPGqA3Qi3fE5ezNJpJYGaCtZINA4DC1vqGriGmu9
FoZHHU/8oJoanv/sMc578v7UdPN+vmrBsggI7Y8rYbk0U3yyHQxAlaztRNdkNCqIEB6Ipkg2YtbG
KvrlTHlukahbyobKavjqe6qYsYyiED78+8lS8TlNtpKqKTvxxsd167apVJXNkRxow3vPrH+XYFAs
lBvgN+7OZEn3aI3RG7fZKUc4nyu6PinvHFdYRiM2+Tg1YXmyO1p+si+vI/yGlgMvOxroXgxsOiEf
n++LWzeP2RK/tDAuZ/9CKqb/Zl7Q8owCPxIiJIWKlSJ8WHKmsKCjE6Vv1zvLVvhg7dXxqmCR9WFy
PuyfDMg5WGbw4KRZNpCuzGx3KOc44l/bkmQ+x7JJcFMfli2Dkfv3xWpqIa1fv3tQjblQ1T1MZT+O
tBKOJ7b9lTbisASNMh0uFWCn70jF/zNdF2udraWROJilkuuL0Oja3ul03grxnmdBwU+F/E4xToZO
b86SVU/I2t3T41SW3YTygv4lZtOZgVcYIPz2S8DKNR8l5JLLiimg41oaAVKZKwylqxQIYYMIJ/43
Af8ZiwUGsTOhrX2oy2C5PdsuMpCO5BNpgBr71WjpuhiPLM9xbHBl5bjcaQ5ql+9GwWhDTK4FRvaS
PdbNZzef3DGOmXqzDlpWD3c/5YJHDvhRlP9KcIeftH1zIm0/TmxVhYV9gaZZ7IdKOUabTWVz7Rrx
uxb+IgNKGMavjixNnmqf6RVv3PUNkrwiVXwABPKj8USeJ4y+p94tm/g4q3Zp1LweJAZKi91TZv9R
hGsL9LB83BGGmLTJEbpDtY/WiwZ/gPf+VBShzG9auwv4rhkuvJjfq9XgeLUbWO3yHvSBkKcGqb7x
Cm4zXUq+7hQDBOubWueT3AstRJAHiIQh9offfPR7DmbFVNvfs/O3S+AxSGJoNaAOWRU9Xx22bSaT
SLTOENumwXfJI/uEPnicC6a60aX00eIKvtmZWy6qk9Ma63pMd+srrpNbMsPE83bbapyoDb9Ti1ef
oD+bFyrOE/s5J4h9fAdKDzl3rfhyCBKWj+F4PNe9rY+1QpoGlLyImBcHuVCUoTEpS+Zaw7NEGefj
xaPSJV2lH4MU1EgZ6i9d0VPROSolfZ+JH5xNT00AEIyCKv9rFTmShTG8j051wHTL1d/EIEVxKHre
1C6YzmdTCv4tqaJrik0z9xknwy5d7bzE+r6qJ+Gl0b7t0OBMHXy2ScI0PX4yZBKLIrX04ix3J8ZH
rqOu2BHrUZQibnP7bi8l6R3RiJJoqOLt3qFXARNSUFi6sxN1PPSk4GTQC93ewsF9AOLuEXJRlOhv
yjTlCDr4iAztOH61Rv7jgVIf3SSKelRevNnyoPrUGAYVa1UsnY+fthlbgki1IJWUrDNcKeAkmZmj
WnsU9cUQ2X7bnabRdTuCISCKOMiwDj533044B+2VmThx3fC9OK1l75MiHEX0bS4Dgb16Rz6x37op
xEc9JfS0xU07kT/BDt370bynzaeLZkqWdpRxbamYOJEdMsyjVyCpZvDInl9H07mNjgvl8w0hnyou
YZ7VunP3WPrRXOmhInsEfYEPQ2YqJ73c4yxnuEtQB1C4fIVPa8AmQhXPxynPwhc7nF7DOQaVcWJ1
yc872/74PCQF3B0zZw8cloTDJWaJGkL1UTCA14wjLc5j3ITCUVl6PoDbJ/ReBw7/hdRHw1ogvSg+
2unxIsKuG01Uv9ZZyjS705aOK5kBWucr7X/GuqgiXPEkGSXSsYJdW9BgKGdb5fUw75LTDTXvHZrK
oxmz3SroboC6fHKntjwghGwTbGbVQB3VJikEU7j8tddi13YdlYkTe+6GE8O0f3MZZDUzJi2hW1NE
rb0ZqlPb5ziLAyZcFibQlEoCnLF3B2jdP+Wjwv2ZijbqRfOBM5N67mWDdBj4QEQ/j57F9eroSSFT
5L6ewQoDvctIIQTwx356cNucJg0HQvY/EIUt4rwi+WyChPBAc6zj+5JTTwFJs5cQkxSGRHOpQUwA
obBi5zPDUXhB2CJkXV/156/9GyNlqZxcboF1kx/f7AZPIqvQcTKiDzCnG/EeMSfTYDMfJgcjB9WF
UaWtwY8rXP2d2iDTDxMiDmrj4rYMztRGBIoXh6HZHZzSeubAJrJkr55cxfsHSBeEK1AsRkSkso1t
ZqxUjp5n7PuK29jpUQnmHr5+ck9+9/v7E+5l4oLI8f2bF5vRa7A9ZpRShMqSeLyMMtNo1uLiab6e
smXknaGmhH5FQ+fLsYmL3iR0Kz3y5Lb3ae7XEGQtZiHEgsYt7/jM7A7bsVTCivrLZUP+XTboAb6T
uVLZ59GhmlcIfmYM+w9AsTBCZQkaAyjdDu5zFYitAmE5GLJJ0FcX8mgPupKUAk3L7OgsBOR8NxkV
FvsR6BKjwgnMmkLrPNbAcS1/mkTf5C5xO0AtCEpSFfJtNnHsZvDgvDVSb8w6BsKXe2nxbvlWo2WL
+dMtYMV5BTiEnmLPvCWQP394bVxD8X0bV9lkpxhFyqvg4fERT+3chnM60GUQxUntwOtrbR24InFN
bGJl2UCHd59Ou15jXygvn3qyB1Xj/oOD5P+ZypfJ5nzxmwMpflryiamxnpxNfBpRlqgQJfCxQjRv
9zcx1a5vypYS1FtcDf5zz8BUNJcry3b+BOaQrb243Bzj466aCoCPpOc0+SHVVIzKXUSEkOu82n/X
Jj/ljJCk+gK4tRP+rimyU/VJCCOoygbGpSoBkf/Qf++wQFGkxSCyroV1p3CeWMkAXmbLAYYv1BjR
ho9Wg3Bhg5AKtIW2MSIx1BH/l61AOr2XlmwOu35+KXzvh8bXn0Q07z+gYd+fFtHea4wsyuRU0W+s
wBG3iUUAIxJe9CcvnfdKSvZbpMdLRJbs+6j6efNH44wLVMJIG4hzfVDlUE0akjwBWj4fFTRxQk49
NM6u6F5G03lXDYjTrtmXiKa00uCpb3P69zt8lWMfdLw/6d7mMC9OQkQv+zdzQp14nfPgIF3oH0TR
e9hFQKKYJleBccGav4Oa5katf0+aAoJOIeoQ9H9nZdyNo/PYh6nVGpHe/aFVpsrwcSSIDz2dr6W2
ordj87gMNZCqzTJrsv7K6P3Ye3QqFRc3ARTmwOROKuX9gE8Z4YzGtYr7Gu8UE8BUCEuCPJN9GEJC
GigchjDUSSPyQK7LE9UyVl3ErETkTQ1GCdjbYiy79HiwIqM3cps4yhNsMafDF/SQDTbmFOoPUxqB
/ApniJuj+mPJ1iOIi/n+nAkgRfCCVebZ2V9s0anseXSNP4Ifgoj5xOYXwxYxM+/6Vpc+YQmaKHXW
RuJNsiBpzZ6I9pPW/fpgl8jT8jBAGgORvUrNXAG1GB1OLttHNyGI8tWmu7faqcBNb+SCjJEmSr+m
z47Hxnq7Q5YOG65OJkwKukK2EXKruf0aggtFlOrm8FUZOOznnECzg3EEM4qyw4xUGF5Gr8/ZmxTm
xD44cgwWIb5ZuRe8HMeDeS0OnWUixSZnhSn/+bgOHXax2PUT3vdsozxgH4UKZeEqGew9b5Y23Kr2
OEZyVKZT5AXo2wVi76I0xzVA5sJ95zCprDFlsfxQxZy9O7N9hoq3CD+WXB9RIBaacdLy4P/2X7+M
ENcpYkAkbIqDj9+p9zMJnvKXVedYbE7EWnGVXHp4Wq2U1uYkyTW1K1esv8DIg7LluynBf0pXyKyq
0UI+ZfUTYcija8Ga3nVR0U1DMegHZTjYFxFJn0D2a3hdSP7sMLEghjbWPuEfS+u66j6sv6FF+PHS
eoRo1w7T05g0t4fGAwmFQZ70HXFC05Ij/muN6S7nF6MB2JTZlmiwJUUvA5uXPj2xjNJ9tBBYwsOH
Lb11+1aiNpQhCZ8C+Ux0viDhzZ5muLYgdFDy0JDJHgwMPZCo7/fnML6LC1iTWk39e5HuHt6Zeqpt
QWHzccEwNiG62Mg6ekBZtEsIYJ1Uvx7wyxonrZ2tGAAbj7zbQ7dYSVIsQuYSB8CChgZ9TiEEU90i
Tu5NOx/EQ7id4zW/Rfufrgr0Tx90ByNMAZhw7LRNFPxrkpD8eImQQL6K2RDQcQX2DaIkFqm/cegD
n9Xno+wBSOLWj7Kdg8AcBDtGc8wqUf7mwymwLvkyQtn+yqu4cUzHwT5LgwD9BUqlPkW/i4bwUlcD
Ki03pRmzXT+ip0j8bdsO00cko5id+PWrKweyBzhLcm4gQ4YojqXyxuA3ytjEwuKabThnqUfb99p7
fAHaYmzIQjIVcNaLSktoJi9oU+G7SdlBThrIgOiVTwlHQEQhCW0tzP0qPxRcZVbZuXqYevGgqEfk
KVbV7dB+TUqmsNsjFJ+LUTUvZakOEP2Acqub0OtnOBB2H/avskfl9p1EztxFrcNviSWTS1oYzzqO
68YkTFwoGGXOXFJWam+c8/4uReWkYQPWeheTXzUE//uFtv36+ZNe6uijW1hYRwUivuEV6+yl1KNu
wq2lfvifSRoQoQTKXcGzHkFrfqovPfWiozjQDlPRIx/nEGgTMMW1AfJkRq1aPoDL5QI//YMMhE/O
darqxQZoyimRKl63fTrbMQC+uwsPdjCnPRtHFSxiUZEaE+sAwd9eAzaGksbl4ks5Sli+4HiSTgvp
xd5obI6Klk0WyrnK1Mg4vBG5CebShTB605kHVuX+i9POpz+FgwCCrgR4OrgV46GciIp5wGfylB9P
DXHxSAYQtvn4WV6TGIHkU9BwOfGKjWAK3ou4XVprx+9IAem0ocp0lb7SfxpX/wVcE9nmEw+NjbFp
PDSe+vtgLVUIhKdF5+4YbVH14pGd5c43OLt7yQIMrVp9kKDMXbW+YcOlC2HpWSAMQz36W3T3WeoG
yhr5FiphPFFa8owGVIJLVd/VJu7BlN9K+xpS12BpZG7IJgk2pq9QD0ftABAW45XrlwpHIbmFrECU
PgiW7QX31kKlFBhiNyub3ejAELsd7RJKC0SrqCtGGXqyb4tl6Em7B4yOrUFGlnhOAhQTpEelDbHw
wVV6NsZBuUSFQuf9heV1Zw2fMX0r6ZKkxm6eCxazs2VZqv4H5u27tu/GD4vXSUCPFizHD8e9uV+O
o3CO5hUiPUJUXyGGE0XqadzeLM2TBOW25AeXfh521mW+xg+oIGj+wcpGYfA14kFgokk2XIEC8PY3
M1rAlILEIS/SPBq86jXe7NSqeWb1zGtaheln9ZFVHKNWJXLx82cUPF4iv84SEg5ouf+HJeQkyQaW
DJExMe7Ihbvqtk7UWiM2uRP4/8je0qxWwhvuTAVNYDB8pH3R45IbCN868G7jTrr91hxpqlcKOTU3
+MUiu2NswYL+tvEfh0UFQ0ovec2jCRarQLlaoVvrc0R5mS/2uWaj97BhY4n2tC/brLHzS+9asd/K
WcNPSeJoGQR/1MSGUNj9jEL+OGH7B8PVTAYMcXnSih/UBo2mu+JcXaR7UOf3+yqmtJWcH2CeOuQv
hmL+gh8IAzQNjCpOSfKH580bYqi6LAYK7h0iapk9w67mm9iSYzCUJZpP0UH0lFiG/sdxXtWuO934
Zt0UaoGSfilJ+ASTsWD8LwLe5yLHJ7DiXP2bukFgjYXdhV0kcPP6ZrmYnmSpBgEPMGkUsKd1VVoG
mXDrRY+gMx/jrgkDuVCCGrc0wmfA0dWhTwX9Z6VTXEs5kT9kdDvxohwSyLlcobEnuuI8vCTFygP5
IN7SWwt4P0+X40YGUG2Fw5t+Ji6OTznbvRbBz03CJHW+9+TT0x649aB3lBIZ64PrYBrMPiuXeYYO
KZrxnIIjmwSdogFlZqjVyxBjRVMI+bARs0l1lO2piYbYkcx7mdgl9WJ98Pvl9QCGT1qAzpNB3jdM
5wGQuxEUFoZdj7S+NumkKSbFxJn3CtOqkrtthj1gEO8UMW3322J996X+tbXEA21RU8B/A6zdd3By
AnbGTZXs7+YIP381YKxONQ75/SfsW30OitXAUMXrWNhyriia2mJk3pyWUmqtjtqrlFz/pQZgEXmO
u/0HH6PHAsQwC08qpH5YZ3WtFZwLlZYlN1XdWfBJfBemwOd8VCb7eQnKwv1zq71xrhbFjMOza8md
fbjIRNQX6wIB5fmHql5sJpB6cYhUuYyZkfjp7w9o3sSovAY/t4Ta4AmmgsYTYU1kStAXcWL4g11/
LMUDPQ7AwulrvYg4B/3kRGUyD6tnq+6P4P2vD5+vlqXSlM0urO4d+ErWUc6y0o8+UmtQmVcHhrTZ
qfr3VEtVTFVxqo+jyTthXu+1shRq2JRHZYnohDaxop+rHvblpghkynC+bPSHKE45UukJk4PW1Jwb
xmGyGRBzmmG3h7cmVji20Pj9TtYDYqqWSCblz/jr8k91gDhqxCYZMhZ+IsfBU0w6pd/1A8oat0hG
by1YSswDT1RNxjMpAFkCDGQU/qBfXY5wSJOKDQDkSuQe4UeSIDGzFJfrZqJIhG4Lte5dsZ7Rv1At
ehpS62OSSk14JcPBma4xa3pMspp66IZ3Q6k5kRY3lZ6KwqHYcNLM4OT53+PffOHb43DiJJeXog81
HPLk3RxvUvs1fBswAWdKOOC+eadS4VHoNtIjvkh0Lrl1pNixTNB+2OWrcue3xLkrSil6ybUImXI2
lv58vyMrssRHymjS6iefkp83slcCjPNvf1/LGEeoepDiGkuG+iZLBMvhREber3iXjLtVAV0WhcO6
Z3xhB8PWRLmqD8x6LV3/ZBvqSxHe6DfSJ1QjX89LOYsX32jA7GE6VT21jhEfO3VJnXTRrmjtGG29
0wX+Uq82UkkpC2gMObNIHe/S+n+8zGbzFXS5AuFmjfxvhnZ5TktcEzotABXxeSk+O3E+yifQOEOa
pW/27+QAlnJafSJ+fehy/vwCv6cobNRSLLbW7OIC9Zyf4SBkTPxbSUMEpBX+BUHh/Fu2Z/GHsnfc
JPCnUWGMfO9qMYlmUZxluOTC41Ecz8vcnoXTdDBSibkQkEY5h49wKIbADd8LEf5eETL6Zh9yvWMn
mao+IAtf/o5wbsmleKWZ9amHWbAc4XtsFFzrgyji6OXXh3nE5BTvNGao1mR45jGO1VvG2yQQwzGz
r3rayvfE6ZMk9gMB8u88WKkPylqqX7WwyOpybJWrKlYy7RmG7+1ErHww4b4uNeNKE8A+MRn7hxM1
mAtY60/CsIsO5nDBgZiFVQkVK4eGBeEgdGdPQjwgc5dFn+vti3ACVQyLOLhFT2ykFF6EH8E+j4br
W8QnlbkrKz53XYUoCy274AHu7N48I20ALI4y+QWKCQtpwdU10dTg9lESzGPZy0mWUo04lOQKiM+Y
wcit1V7uRFy5hVGTC4WyNlLzr7Gz49KK3OG7CUvYj96L0szEqVHsad/yULYrSSQBIUZVjoyPl6QN
VSmvI1O3E3B4B/kYOoGQsnE9X4zZSFPvSsdcn7qynjsIajOqtDHMt97pwNNkD31D02mAbM5gbr1I
BmPT3Rrm3vpGoNuAT65x/SNvRfDbffyZKqy3pg1hdXesAM4IAiBOX69xCY5lTZj9CAPWqEhGzbL6
z5cYgcSvM0/CXkafxJ0cj2UlfTdhCxoymfJ7f108u1i5Sce4TTF7Cqto5pMVsl4bMgtzfCzpkbQC
vOqePIWEBz30OLZd+mau9esFlvhQ9zK9molsLgvW7AYg1NjBQm1PRXPnUtFbLWUCl5uVOBJc2qaK
OJQckfW5AP59UgDGDrzwv1RHyGbZ9JC2vDiPGVvnEUIuORxG0MSxPXQZuuiQ97MAG0VWsn41MFz/
IKPnpbutiVY9riVl7chRGO0mZkc/KSXLK4KydmBaxV3YRX3x81ctdLRYKZDDSZUxKkei289dENLr
qGqmIBlvv6cLbV3p2OMspuiOqaF2zOk7bR5fVOpPfiCiw1IK5OMdvEP1W6VQaP2vRuoIVsFwzJJF
SdfX8wi/b2Jpq/f2iBAQw99zyRAqJwbY6yGMrx6kcjLsPDpPuRg+0C2orM5WJ1dB4a7pxHD/iTSs
ULzk0+S8uG/dSnk9FGFWFoVL6ZTF5nlD4Agm3iue0fXl1qoNY6XrBZyqb9iUGl7cFZNwhA0W9gq+
P4M00RONnPWmFlQwmXz9ZcHbIEZVU7ZuHFxr7yhD4OjVPoghsF+UeVtQ/0fdsGqn1ESBuE/Ro+G7
AFJb2LJ8P6Z7tDZsc8hjHcXUjufKY5xv53e00mz2eNpoUunP4eX9JgDVLJY9GFZ//I6iIna4LWIS
2DkeBuPvBxP+XOeFJcM2spH1t1IEruZHQ3JYiYA4wpC1KNmpgJ/ohmYyBtBGs97AqaL5ArOoJT7y
jh36E1gqT0wfmSG4Qjfo6vXAjiaVRlkkoJuaOkd07vxPv9kiCn3xvKXlnleZ9Rp0WoUVzipDJ6+O
umXz214M3mRB9JZlMKkXIUijdSuWuMX+uxKZY+mROZGqaZjpvPaRsKZHly1SPRBLQ6LRXRLqWHj/
1S0I2naSR2oVK4gslojl9qw0YJPVV2yVNmm9oJEkBeSTpjWHqC1e6WFUXPsd6/LlDs6aJtmBdDDW
qLWxvR8olbwqGOwODOfGaGKfnBgM+NgwlSse3lS2B+6s0Pltwel/9x/UWSdK882Ecqi+bckmL0U8
IaQTFI/fFePtwEJ7PVJYrQmohUHQ5us6eN7+on8oTnO/TQK2HkvEMSQbltbOkaOc3Kd8G4EMtyJf
Jeps5sVlMEj9xEVh7o3B17b2yMrnF5W7fwLakBJFtlbkNCbOoKFmzbFui/pY7DhGenuV9UYbX69d
k9EGR9zusGimisSxl9rrJy1a0gpLr0TezDAeNgbZJyWfEvq+5V955n8ThNHvW3MaBWZ5bmLKhXpb
Iq8wGXxriLvHEEXfSB0oTFffmW0Js4w3SprvbqN3VSNOCt4ufiEk2ZlIrYqBUDAFWKMta6jzzf70
QsyIcKK2p99EET9ZKCYxNDnnCjYwQRH5ksZF14FtZZHv/10bdISPVWEgBd+1Rv5PswlP3HJhWFUt
zn3MwYediLuUMnPzNgyhdSj3n+PgX08HHYOpKGwbZcPNbSuSEvrebrj1reabSQHGhhGA20WySJjH
RlHvSe+kzjjI/Y7JnauzVUt7x3y3C6kuFSzZuOkYfdgxMHP0PLx88NBEC9gws2f7GPqXkLrmbFyh
GmguLKvvV4go0JFXhRKzlVTrA0Sglew2+mtm2owviS+Hx0x9dH0WIS12520k3jnK+XeawLRzKwuA
O2qTIJUH0AX6wLXljyp5QaXfbXeZp2szO5jj2x/Qf+9R5SSxjAKH+KzvU8T5Em7Man9TRr1HyyP5
dVvufU7MdPGtpcMl+tn604tISG+spSovb5umBxIl36p0Fvf6jMf5AbKZ+p5+a8B+uNPhFAH8ST4U
pwEg6raq7nYp0YoZsiGWU7q6+cM0VzI6ZmZtCK2Eq+lkF/Bh2JML6WuLErFxPxHhYF3qjypnikqi
D/0+vz1mvE1W0OqYYVbuWT0IvdSLOlILSU/8TUig21/Q7I9DJbYx6p7OxhrQVumqSTK9JLl9SgoL
fZiG9FYSqPRm3K9myVTg5KOoFSwhkSzjisDko7w8KYwvLury90wuJhv5ka/Nj5Rwkb6dYUnb1xNC
hDtDW2ZEdsmEMge9SpUAB5jpq1RY5XLurX0bWGi7WoO2WXk/eONHYNyywM4nRL7VAwjFskhwERyk
LTZHN13mojMHIbshzfRHeeGklGZFY4w7+NZYMJqaJcfT00Rdj2NvKh90BFyYvkqejzjNPbHW887Z
z2ZxThKAAT6oIWfbkfTpL4/sQehmUDYqGhmtRQTILZ2qsoPuYTWrGrEcDqrsoazcokzWeXLinELS
/Ia9evNqKy+knvNVJpBD1ur32DQLODpaoHsXJ/ZZbkHPqamHshfzR27JLd+BdUmlz82EPQ3Ct4MY
Z2REnfZRIri1Sh937iz3yJzo6pDhtVaBatBL9bEHCDmkKobjSDIWyrraoMGJmWTWeMnLx+Rjbxju
9xdIdPnfVE5EQAMQMYfommPMh26CEILuTIrpPhYx+cp80KU6ko+cwIA7WtrIwPtQvup/mUU2RiKM
lQbzHBt1rifT1dbx5rQLT/T3iNW9JygX7k8oxhnHneXySDW15YtvpAovdMT0/I1WECaPpOXrBvQ9
zR5uAyFo7FG4FfB5wC2jrlSYqibKDPIh99fxQbC75eAZfNtY+xAXSat/LKKghKxIWfqWa+3pYb+n
2mjI2MAn5S2forRTBhSMov6O75LSr4M8yB8Jab/zjm2m6bAoGF+ZQgUmI/qhFRGj+CkVAJvEGBWe
T1tlpPf4ZwrF7vsrwlIyVCifWZLwMTtuccQxwlO9WUb5ACc3m3923/dSXLjAAfalDqSOpdz3qERN
3pQfSgGyfn20H+fg1FDZNRpcZem/q+f854I2FHUUF6pjfXf15IlOcXNNtEKBd0+7lyYKjECtu2Vy
zfCSb47vpHzOzHUmimcOAVl1NqFMzbXrctCne4jc0v6lwJfEsfoIHfN520xBNVKEPgkVyKwI37Ud
a8vFWZjuLjORHj2GU1O6IRd7jMgult88IZ3nYtBHg5gTXZ1sqII0YkJBNaEkCKkKrq6amPiuTtI3
hj4SI0mfbSnm/z/uvlpoghDMmKXTmMwKROSVNwwqTvJ92g9+DWT52iMS9PDRrUfffX8iGOIkgGqZ
mzYjjUBmOtg2BF59WMPv8OEiMPQhT786PUBMtCFOfx36FwoJ9T49t/qom42+MHMW1BpEQaqRnSEj
NvQkudXv5lHZXSXKpB5qhGNoXCaih9fohR3ck3T5mAWqUAV72DkIX0HqiG9Kx7TgX6RtBqOz25Ce
55nSF0jNikOR5iDWsmQX9D9R7iL1uT06uzit6OOwRvU+m6+GNqZvKBQ70Krzf1umt8YB38cyZLc6
J34L9zZQ5AJHmDPJIDRt8OhJNYqnsTcd6+veTTHZYQzt8xQxBn9Nd6enm3j4H2Z8gKe2AIuYH/Xs
dqG+1e7hYrlmanEcIB6Ief9UkrHUfN2Fg41iG0/rPokZLH6ktoecJaGrrKyysiPsdyV33Da3lpxH
tGOjQ4UfWwGI3mbwcRmsfaZPLCfiC/JM3Hk9KooxbODw1cbTSIAgb+5G8a0gdoJbHzV/Fx6NPqLa
PCVj5qVRPJQsg6XOEyvn05/27rTKfTBAamAjhVOZgmC7Swm/7dQfLyr8OBPNCb6uB6CRbcFFxW5H
MN9f3zTD3YoOEQ99r1Lst770VRem95kGK8O5TMHHhT+/sYg7ecWa6IIZQD+Yqla9p2g2HIt0khOo
aq8davFUHsN6SksBJNuIF9Nuzju+4wPiVUDB3lYEqshu/oNRUsmZA4KB3eUh6yYq3ooLaGvacxDd
h2uBO331DGgDLEzxo8cfU/jwJJ6mXIHsYaoQffGG2+oaToubD6IdZJL4v/KGX0+7MYpLhxX2nFPQ
2gq7/32dfqTw5njZ6oCLkNPCq3KnDCnF2pynUBuyiVgQx3WL/87DWg1anUGoUkDMYK7dsDfOaZ4I
q/TDySKnsUcVdboTS+uqnF1lhD3Ky6jRbEIz4T+ksiS11jgxh8aMFqymU/lcXEKo4APzl5WB97Yq
ZqG7sTvTdccL8yYhL6yrSDzDJ3Xiiq/siW0M3izf1wBxoVUqPIP4VbSu/O/e5UKz3gMAE2Y1b/XE
Gmr57DyTZ/GeDqtfCMe7l7dg+CT8B80ZMWzL3UH9ZNk7ZAZvIrzW6bzBdQ5K17bQxfUc9c4JvS34
v1G1jzFttmncTB2zN1DKg6MrFj2MUsY01Q+Zw2lY1Y7T/ZbqEfDFrbvajchNgKX1YhBrS7toD+Wf
0MVgypSyLmEf+CIuwWMbFynwa04uAnMdnoHvssLHGBffFv3SUv1QzE4L0PZCLoTkkdYoGsRK6vXw
qmGWH8QAYUDgMpd6251HY5twe/krpQM+vMtM1eyoAQrBh/yVl6879he2RWzIZqI/rV9tAwdl1hk2
Fr0jdyN42Yn7o06LENzk9EMsvsgwCO+UOvkmBbdIyGZyuIFg7NljrN8T+aswWi4tSS8aPQFQ32If
Hfs2PbDFLSW4aOo80AycJM0Kq6uz9d80B9ge6tDZRyNsAGCnGI1NqFbWL+U7MZXRT/hifIX1LlYb
1+DfcUe10d03PwV4vrzIcMlN/PVMdbusgovzCtPkYDXVmMckgkAXtdZxwNrOa+locqQbS0NRdpRC
08qvZtK2j7cgjSepzpA9aoSWsO8sixPVVgHzFR5E+ceyKznIhRwfPnYP5+NmBhs92whHloFZfxut
/8e3OapQVSRZRVcx3huepMiW4cjZRSuuhKBrsJLK0kaY91GZyjtuJaqNSZzD1eg/G4EFsTWlJzaL
5o5qqIL9RLS6XA15/nDs2zf1x9T6iqa7Lu5G5zcYjxBrg7iZWAXzCfC35HY8acbjmdR4hI8QO9x8
/zeT4pQpsiUKFtQD/r25xsfeTjf7cvfg3H5JUZdBk0KgmhOenBz6M+tud99xJ+xAeS3/cipILo/y
DixB0xzlGn+SvAkjHBXXlu/7ntkm8j/wAfQR6jxQciqFj7/L0uf+goUGIbJXI4EBT2qoRp0zTGD1
noceWlSoDzjVcD5ePnI7LHrWeZrYro6Kt8n4KjmVaG96ESPdiXidBJU2xtVM0+BOtffo/2bvGcLX
BIvVbqLV/T1UP5rXvN9Ce8rySrLx/o31/E+RZs9bnUSQG5n+CDwo0lje5kqzkdelHrUxl6FcmuTF
lvM0EO0wtqnfzQTVzyQ+7dxzRpCoOZgzN6JPjMce0g3q9OXG3sqkP/Kj/ZUmOQ0pPGkXojXZ0Ujb
uCCfzvcFxMAp+RaD8TR/4ogE11cDKFXdd6ICdzyzebcX74MKAKPsyVi/LG7NvwN4CDK/PHZS/TwG
nBBVr9r9BGLGuKqsrdC/k3PfuZ/4lP5Zuqr2EL6IWVWbIyvb7k924RQSSdCkLNtHGjWph024Q53S
atdCGpR+yyPZnceoG3clKtyvEIOdDDCSUsAn0BEHDMS6RCIiC+vJMc8YBUwR9/7besydBUH1o+Yv
AqVi22dLMntlXTKvvOY8d2SnPWF3xazGVUXdhDHXCNZDy1D0QxwssCY4+jtYynA2+wvz/Ek72tRw
IBFpNmLQQa9kP/tw0nE7FFX7iWEO0zczzOg2x1lLoP0adhRAbrYvNDzlPwNS1X7If9KrKOh1HadX
JPQqx8DvSlwDqNdfqemYKkn5yWUdo4mA+5HXUNqkVlei+BZZKwAcEtpdTljoiK5J1dmFbATl4He4
cAa4ksH3oFhOdbftC7VUkm1bVQCIy6AJhRBZjcMvFtOW9InmjaY2oQiJ+XjNElolsyXu+VYItUvT
x4u+PZavY4cYJO2oGSKJMWONFbafZLmngPFuxzNcmaQS7D72xt7WCn0UEgLhR02mtnCRJT/SZ3ls
chzBfX8Fji8Vh2O2TMfh1xFxdMrYyGQlIMd7qSF+C0MFF7zCb/ZLhp3NNenxtYPp1Ye4jCKtczE6
zQE7KMlGaTktaU2nYHaq1w/FFaRbO3SjIwUf+fNy+QgzjfcLUDd0FMuADyoOvKRt6B6FoVK74F+U
Jo3VHIpc/GncYhlD1bKs55x0Rn5TZJ6+5wo2F4ibibnRE8WwI4ylXPnLYdwUVJucD5fEHOkY1Yrg
ttI2N2EOa5TWw8TTWLCRdYsWug0RwmVuTeOPlYK3J7gU9UgGxiyn8aDxDWAd2xU3ViWcPM9SkG+O
DwnxuLAHLXE+AAmMPcdMHMMK6/J7HXK3qlsUW/XTRBqkVd1VRzxdyoHtvPOFAiX8eXSLK0eRgfhT
ZIyJ/fRMj/F9SXRHuhsPp+7VzT5UMdi45igMG0BwEpsjrpaAMfD0zQDJH9RWLCqCkP0hb0RQrG4w
LZB3/W3680/OY1hTHSRUBQbZT11wyi6XKxNrxIV7iibCLVm3xmX9E3HCKiUmS1Hqek5u+Xu64ts4
2cOLXqH3D6rUGvRqfqn26ea2zdj5Y7BEh+SkPU9StXYMdykLQPRugrUol5H/KgoFIQ8uaRqnCC2H
JSPIKiN/w/nUbT9a0sI+W1Yy++zs8A5EvYlKhZq9fMtKCCKy/7DnRKuezr4F6e2rbWmkztq49nV/
mCySo43jYO/rjM2RfHchX7hUwr4mCChePTEWBvoNeFdSPhuqnyKEmgH66TuFObryNM9LIpEGewaS
x/DVKavNKV2KCNwqTZaHf49q76FRE14Yvq5iB9c0dvfQ4R5z4Ig9baWp5oui3uaaup/Rfqgq/vqW
dk192yQOtd64VWm7Uxbmmk/MeRu82vQ+Z2jpaq+Q0LbWBT6rNYyPmUphNrX1NAmSEBLG0IIgsqXj
EN9DzZZWOtR+FG1fCMJQ/AOXCimBPX/UdjLe0bIucNs1Z2yX85Vi8HH/FTYn6BRDRZMV3OfAM4jh
7n1i6mn3NLLqx2/8PPb9Cf7qgXt9U1ltJd5lHZNSDj4DJ8R9GLbj1/kSzCNXnJeKo/WNUzYystlK
zljMkQUdbOm5gTG8JQSaWSnJnNOILOHbzC0R655ENxbXivL1B5WbHsRgU1+5REnXeWRg88BCFln9
fJT3e+Dt0EhsxorveW4wv68Skf7nr36goKDBpa0FKAizXn898tbTyEPmq09jUPfk9oFYyVWHNra9
+CmXnbh3yBkS2jkaC2c7wRu6UxG23lVVoSEa1uldpvqi8kdNFT+1cJOoNr6LHBjmLIMyCfudYn8X
G1qV3YcQLZKXqVMHZ8fZyB91UZZFbOQRS76UF+7h/L1FOpFF0NbySf7axjxoXilsfsa4i0Bw7zaC
EQm8EE3brmJ/mWJwfO48/NZBmZXUKSA11fzGn7zXQyyJKhKaeetXuuBcbhcuhDmI+712jIGf61v3
Hd2m1QCawjb6mJgs9/gPnS+zDTgdIJfqb8l78FPjtXMn05JqBhfAn8vQCDgjd2dCxDd46+qWF2p6
e5LB+i8YLRFZ5yo6iz4lyERWZyBI/zaSlfNblW41/jh7u/a69wnMkW+dWPWFjkCTZei13oX3c/DP
dPIqLoZglqt2W+7PsW6DD+k4cVSEwtSM3onRVNDvUJDpwMde7POc0xKC9LlMlt/2jANyXjpsAFCU
9yCavNrKd8+uPmPVE/PJrZc46sS2BuQpzocHSMuSU98YxfcTRBtMUkAs9fftvBVGk0VJZ97xUlPn
2JxBljWwV5OgIJsSi8MZx1O6NyRfwx6kkb78W/WkOTX+X9MUa8GEbrD2q/z465h/YhFCPqxLrh7J
APGWT8g4qpo5P4cR1/1MBi5X+1lDSqtzkwgMtzHnDG+Njk67ynrZACOCwCJpN0h82E5XCgMRaAjn
0fO4lutR7Gtz1ILTwk7MyDuVU30u3/GTOCZf520Nmbyvrh5Dth1a7USmUIh6FepnSsiDWy/NO3l5
/yBTJf6KHMG4ZLrLKjUnb1+oieebmgBL839xc4O/fEVxDoiQXSW/OktMErSoDqcMrEOsFhM1DTaw
N91jQOR4BcJkx44MBldA4F4zxn3b0OG62De9AyC2mzWzYyStRMiJjbxKsNIHOfQ/G7Gu34iuYZQg
dan1Ul786yA815dzsENO15D241PcrReTt3SBrt7odCc0c6QYB3VY8S1VbgTo3oLROTwKfNrQ8Efm
U9/EsJaA5a4MUuUYs853EJeMkUNu2eSCeMgBgMHQj3aL1dA/P1pJ/SQcbUhOUOClc4QYgmOtcwNZ
6+/OA6Ts6wfAWJqNJ0ne2EFlP5s83ZACvNpS3lqrheEAVB7LoV2AMgbq/cJ7m8zY3GPwwC0XbWPr
t7DpUkr4TRd5A/X/JrJsRsxMkyo07xVl9BNKbv19PisIMjBHcs79jHiUQWu7YrSbUhudoPxa5HqX
KsIpMKn/RY4RNxlqIG+i0SeHfb04TTjeWlXLRkyyI5fDKETL84Zx/q0ONZC6TwOuDgMybOHqtz0R
Yga6PvrtC45e8ydpf+u2MXabyCp+u0epsUFBJVF6pB8YTlEAXFi6JCyX/ILGOfGDNozVe3SA5NRY
AJyWdMe9iCXxq58skoQnp1eNLvGAlgE3beku17xxxoaZ1glqUrpOuholS8bRMZ/SG6LAp93QHvhX
gtyT6cB1+xT1ZiDaGxCHE8qTM066e3QFQ/dXF+L5dYSKjLnNGeYHZ4GXPvRWEwLBO+LKoFGIjd64
GZGP599heDSW7th4dI+4mmJCIkXRu+aGJfYYLHT+M+3R807cNkwDewsCtXZDccQ004nO28QeyQ4l
ZFQOs8T/zNv3PmS25vk/+JALH08EpTG0VrT6htpiQHYIuEcHN2TuqypiT4FFipIl+lVHRszKGmMq
JiahRsN3NqRHHSfx49BOq1kepdepImxEPBLHWkvmbe36qtXPbjV+SRqTCiO/ZpDnQSs6BlSd5xme
BKVH6sTH3tt5aLKpS4vbioQH3Pf7fNaudvpzQhNlFSfxtiLydV6cZVMEhy44nAmb0fVU1IJSQgWl
ltAnGAAxOJ7WVNNWg+2asux5MpYvY1R/4q3NJiCo78z5us+rgOmc6krLsN2S7z56g/VmpxolVVJn
Zu0qv+KijKSVpug5fDrglJHRAEXkYJfWeQedNVS2TbNsw7WgfNmyuDl6/gjx6oFZ67/xMVe70pKM
7654JH5gt6Wh6O+K9RglyCALL9PsLt3sPAwpfLH/C6HXSCcOccaXjhkqbs0m7u/LmUIl1aPtoQqq
ytLW2Uf/xvYa8OnJ+/yfxeZw/IHTfdlTkJfVCyGxgjqNdB4yBOG/uURLHdPMjnc+jlUwWmyV2DB3
eppR5Xn5wkl8hHmBsXDxvlAWcQYgj+POIZJmJJJYXjbQ3AN33SZUOCj4VFj82URAAFDYFcF/m9fe
Omcc5bpfbBDrSJYjzVBvUTy/sLFQgcMxcTj5hZoMJJmw0y3AQIlT2m1Qi429JTMMwK3VyMIF/Pm3
c/JBqwtse8HcDzOziE4eXYzp6rvFiuQJBVDDRcIQe98/jrIc8+C1GbkahRZknMNhusLLf9D3JGJk
JuKes1R5tUjlOsDJdk4QMspPGmw3tQ7PgDXK+qUI8wVEbr4biFLB3VTWshQsX/z3AFGVywVrYp3p
01tprvVEucoyhj+25cn4jaUyzDhhxttgbgHNtq+EXooFvo+0J5r2fqtUJ0Uv+VfU3/8rZK2xKuO2
0r71YCr77Ainkn6TSR/ZJIgCjk6+1YFTbJ/+xs6uwF+6sp/6i80gqM/Ahd1J5IyUwDdzdQsXbqxh
RvUTGz1+avj19BqeQCOuMIbE/NTzmJKEky5IxPOqsqUNShHMexQCkKVjUn7qZyCqEyRD+aynnm8J
D7c19uS6bzTev/44A74UGtq5SEgxNjzaghAplkkkXyiRBtGSP/lxuNBmnHxOVChHsk/0zS8dS8BJ
T2C/mGI30f4SwpDuiR2KyweWEOhRgFao5tDN1XUHtVisdovcxLuk46pBAHmN5XoX4EBO4vnzShLn
kydPnZPgAu35xbtszQv4M/7GAIXYXwGj97PcrPpOaxlwHCX/1LO0+CWSE4L1P1sENmOuZWlGcu9J
8jUF9Dw0lZZREGaAFkd6eE4DoTZKymXQmlFuvGQeQkvHz6WfI0do3OYn50XB062XAAcckpt7NrKh
wnezWq344RiOj4KMkdQB+kx04seFLYsVUU4C0h355KFIHRIoeYAtqKLguCc21O8bn9zipxMKxG3o
IiUTNFFDa7phqW6JqE/mlkarfIjmCLtcp9l+zGGMpNp4BcbaIsgLYxD4X4zhdcOtRla45tmxbevH
N1M6c6t4PF/dnrlagnIAKTy3m20rYLdb+8A2Hb7aof3wP2HTtjDkLeM6a33sVQCNPQ35Bx8U30vH
mEcw8Mn7k3+HaYOGHs96vRPCqqkJn83+XLq4a8CYY/KEyu3XCimZeVr5Z3TmRiuGe8FU7wBwl+DB
3hVkhIPMhalxlngwPbXr/evStVkRN6lHhjVahAFki/vq8NGF2ll0aUm8wGviw+I/HorgMqm7gWQR
YeKLL0qLmlT9cMcTNwOe9yJ3+omWC2MmmMiIWVcNJ1BGJhkoGT1k/WmeYkRYm3Hre1UBn43Knugv
fce2bICXXxMo4t7NRmQ6Kq+xH4zlLqiXNO9hNuGgAg97FjRSi67+dW7a3s8MKQbaZav0DALzq1nK
S/4CmxIA+7CsO33FyGQlAczJkIq0aDQwfOKXvAFEcy3Jo5Dol30EKwtGvfUJWNraO8lqJu4f2z3d
VBhAa3udfqGDrfUt4Tr+OYdbgzUCzn3ZFhepEq7SPCZtTCP1hrCjVclsJSkTsK/cdsnpJrCSPKuP
mvkXXft0jgi91T2+h6WYglHkk8CX3MgnginxoWcLN0x0heDVZHSfozTfrr5Ek3U/NVA/3cQbD7BK
r4/2BF6V1pum+zcgFZhNj/ILQ0Rb9dq3BgbGQN+LChXXd/mAfwGCAvYxF9AaNXLBaWNRiFR7buc7
OuLLYxpNNOyJ4Tb7bRnFuP7KCKKHhVeoe1ZZppBHN+29+e/C1EfclJJcFlUPGSB/n+WtLpcZkKY5
F3/HWQo+ENZCW8Dd01aM3XQT3yeYgMWzshEkF9ivyICOQo0zo+UCS5F10iSqI1+baU9Wkrlq7yzf
nkW9tgbarDH5isoT81SsWY4m072tDsoZJsNcuBw/tWoxYFRfZeRndtJWIh5oRdMrO7CuZkHVEBwg
wutZiNk4wHdSzXtQwHGNm7oISSFgLDZgttgY46vDGnGsNpI3MfxqnAr1xl4Gh+EFaISymSojKJWU
7cccOSHjCZ+Yw6gw2pkSf2S8TuX0TlNMKqR0WwsZsEtDhJm5Leq2DmbeLf1RQHGKlgoPKTeNbPFu
hTpuALTEcj1GEJXWIesBlQ8nimVJgd7qeQcnHWqPNcY9xck796V2VvZogadT7wnWwvHUmo98TdRi
oKnU2onH9XGeG9wZ9s0XYhJXDrVVjmYJOnWuCT+pBW+qGfaEUVGTIhmx0+hzrnmwik9EWSjLDRPv
CShbJevkfGP/1lmOFcqFEvBcbE+1nY7YAHw2mdzzaXm3cGWzjSYPPLdPxxeEeOkvCimfRFzl3qTj
/1Z4U7idQ96+KjLJMopki+y3B55ChjEQjN6LQY3gL2PRxf6QikWSZBKGhL67gMrhjUt0HtUmwuVX
e9OB3L6Mrl+1p8jRoa/WUdhWwz0g2AUhcmtWDIdjx9WveCdDpfGdir8m/zac48voB2ZHUFZuCzne
5yyXhig8iroTsCZPrhb00BqnUgolkm0ECc4lru6dwQBffIwO/74huM3Q81OZw4Rz2+5NLV7+LXty
aeQB2sOXZ13dCDxvu928r57iNeVdmnvMjA0QJFZFuKahsS0pDY5DGPrV2X9SrZG+r5P6v9b4YLDD
D7cvqeNl4NkFH6ZdcuPyqmCg3X6LMZHarX1fBwJTZ2kI5IkXW83OM6AejXH/RY1ZtWxdMJbad4I4
R/j0TUiGa6EGBQwOF6KCMRtJ4GwMq6HHhYI43NQsDETvNSKW7kVyN2kB5SMSU/gHlgeQKoQFvhZe
knLKb4nlsYy3VIEUMQ3yR5pdOMyPkbEGj9Tamvs0HVpjjV9n4YQCG1SsfeX07V9+Clu78ktXXlgb
TFuOgTdtcNskn7pYRwFa/sXx0p4hJ3VQUyW3xEiexrKBvqALQajS/2ie1kHzM5f+P8BnXpQmZaPJ
A/1Z3tHaw0cotn5BQsibmB9Jov4LpYkdrBshIGt1bUMyzFXim8HpEmm/Xv2VGRVF+cSiGMcrpLFI
Mvxz0pGvH6eeCeZZl4MXNcFWQoXS9LAjl8Tq0VndiRwgpH/k+L/0XhozVjmTuvBvQVPGpuKcXYxf
64ZiBXjEF9gMJVz/Sb5Ql0Lmu5h7ChJrMXX5xcrgTqybDStMe7Qg7LYk56JOxGlsyzv287OiuXzW
B6SZZoRIQ73G0UwN+0fT5LmlwDfnHWbookZ3no2IjXfqVFqmZ5e+X1jXoUTwLsoL7+QBSQQw57un
ozV5C2IlxwZk2ixPoOeyaPuw8/qoGOUjg9YORve/0TKrTt7WtounPRsz1kOiREdgIazfiNA6YU//
9RqJxuNT+zJvFVbgJaJprI7vVPyiqEV32jpDKouAH2ytva5LcVATCYPnI37/OxPZTeRL+fsXfIly
Nm1ApYyn1fSZSfuHWenP2BwZxKU5s9mGyuijn7QA4oJAwwqwmwIl0J8SmaS8jRAGIEr+wJLzYfLA
SAgeksHHcu8hMoxhPonkNo0Y9sg1CJ/hwxN5Ei7FWqO7HfR2zWvZKA95QV1r/55eTUSjjJKIFk/w
iLNVEEJ0dkaaBj+eZhGbNBrHC8MEt2RtrmHRTU+LNxv3juYc3Z/n/S45RqQ6Mklf4zHWGfOL+vP5
aW/qJ7m4uk2wxg0uo5oznWAWK0dzdnheXpNSpEOuyGSEeiKPCsTnvNKJJZanZbEtIkQC5UPCuOHH
hStcUTMdyI9URqjdEnSbks+ktMuXvm2mGSPh8SUrc7veFUWXTdkRPzkneXwDo+EDySSC2ruH2p1z
LBg5xgnAQ3cfw31T0H1fXYX7BLadvTGQjfV2/ydsuE3A1N4y2FbgZ8/vr6OCjCXv2TG+Rn+AEp0Y
NT63TnhTpX+1vl5AZrqs0V1qHYI3tKZJdHBut3DT0rV9Lvf4Yv7f7qxvaFKO/Q85nI86Ukk+uF2v
AN9NatlIKe5QSRSXJa9LkMnDtZn3b4bDwWhLpycXkdrbjlqn9fUfvzHEBp07w7KroWLhVIbFC6gC
qRtmbBgBhbvYpTR4kAjFpIPVBvKJwcy8kryR6B+OIbxu0PQ4TVrQLwN2L5x23V0XhB68L0ShjYDV
dy+vjuX0DnNBVJfYX7WYDU/VkwquWvgxM45lG2K+UjueS252M5kdNy1Pg6XBlJ5mqYktfEwJHT6E
+PzFEF1Lxfypzv9SNVdgqHdthwdB3sZb1NRy4IUVgRAPFi2zAkXQJGZXvBVg9Ij1OYrYxC/P6TRP
D/E9GcDssz3/Ksu8pJ1CGxeUSP64VyPIEdYzk3n9o7rXctuov9DpHZS4MzylBKga4At3Xvab6vp4
M0v5F2IZwf3yHele7vB8UjdX90Fbt5DU40d6CYB1kcI5BeaextfibkE0cDyC3hZYqKGRoxYeXgGW
j7KEXLi2pYcwgY3pqvtAs1dyMHcHDVpr8imxCT3xZoLLle6YnyuSeuBXRP4JV5gpCf1v5WQkbyuo
PTSWVx3WyIf9w5T0pW3vtNXXI4nzn3j3uBMiXRnBQiWOcsgPRdS/TY1RqKtZOOSZxDWhBqPpjgVi
zIkq1dQNRt5Etx04zmuP0Z5MPYQD/zAwYhHjWCUzwwHykEeh+f/E2Qshb++zKxdpCnVPbEPkBTgJ
ed6C+EAljVuD4BuXZfkA+xq9eL3mo7HErXMyvvHAnGV7bzbmg/HI+TO5SYqBoC40vQmwHPcyPTM3
abu1JRjTd+aqa0auo3OL0NJ2X0nZhFoyssXMwiv5wiPdgUTsvgg+Y6GgHKz2hXtfuA9sULjlw1M1
2Dqqnkl9zh9ZwvwnnskTN2Vo5dIoJDLAVCstIpSEmvey3geF3s2OCqy3FwC6672nZtMuZRXZIt7A
IyjPfBIKdXNC1YLDHpheaQyu6VHYLGYd5A+HCPlvG+XX8+UGBbCkVyWtGt+LN5FDccSAlr3NEMdv
ejFh0bko46CUQZYLp0lCJc1zWR/zUvPXOeKYIYV22tFWK67fgITZ0rR4GLyHWNJcfpVkM8ALXGEG
y1xmRY1YfLeD4umDHEwBKZO64owI3Oy05nCwjjAdJa1ArVtC60EAGfbPaPGE3vcGvhc3OUKGxG8v
0ew3gbsj+unNlW4N6Re/gTQXT2pJdBqxCLvQLHu+cSvgTZK4vKbhBu8ZNsoLeH2CCCSa+DMz/9YO
KeUbSTUrnM24e8xogfD993s8RxjQT40qwIq4y+TGYC86f090raYTv4w5SLSnTzmJxEYn6WmY/67H
GV1Sn9++LlfuoGfK3aJHej0TV9JW9BzTdaM/yG9Z/UIv2HQe2tlqnQHB8gI8lZMfB7v723Y+D0iA
Wd0yFqi0X6Ma8TPx5zgx2lXve/JC+pluS3D4BlZrqWrlbXzZGW9HynztbuojqmpLaRVh6QWjseVM
9MUju6Ckf0tJSGnx0ZMohcDGziGn6FxZOagvU8I0hwYN1s3/Cu0OrcShvHYisHKMTY/NCn1xDbeX
YsCkADVI5WT5ZskVob3npnmfVMcG4uL1S0uSh5ubQ1HjinKfuK+UOYZWPIcvdtm/s+yX9r379Ioz
1MBoYo/tWtgHxrOXevRKsLXjBGEs732U9QQBDbvPvEeCDwjsOw3/kzhH5Lgi3ebuiHlySS7543QN
JhggY/84SQV3bRKurXZXk3UgxM8irSWgcneBNpDLoORghp/880rlCS6bd9NlVwATudP3kJH2++y+
ZB8V2Ou3StldfM1EJPsaSioW8yVxZuk4TIswQQej1UBWzPZ7SgmHw8EZuJmM79Ml4et9aPSDjnc/
Nd8pwhHJUX/lX6aGZ9m/eps5fnkLsSmothybqgffhBvblc5T0DvV4E5yDU3WYA0JS9DxWAhGsljT
xvwppPKeyNRl9pzRualp8g9p+RMdGajx1CajgPqhx9PF6u3nsPbeWVtGkpv1r1Zp2x3WeWa9tMVm
T6eVPlmH+jW2hsdl48+GR6jzPYge875LARncDE7Cg4XI/PqBLdKOPtpdQbif22eX5g2WbTPAApNr
TVgjFXkMUuyo0h67zj7raV9t0DtGvWAzA6h6PGMF1yOvFlZapFk9qjj3kUOnC1VhYNsRcbFx8pJp
vUemYBUObpS/saGCMBfTQowoL1Uwinmv/ReOR3TL4aGXTI/cqzO3563Re0fFWnQzIIHP0YOeBANA
QxlRO7xqg6A2U9RiJP/qCfZcWSfXiPIeWt93hAK8pm4MIEUpX/eQvZu1PN84m5EU+tJV95C3RowR
mVxAhiq6Rm6Dqp9t8ME1weFn1X4/KihAjsenAD/k5qL4AfQm9VjZ6BnONimACZ4boWiA8O5NUoX0
NyyCQLPJcOlXIXsP7lt6RJyj4V8S7vOyqkF7Ry2yKDSn4XxtDxUU+NS7Rhv9XZNWuM07vYNwxJsE
9nXdo8arin9dmSVk15z5ZN9ruB76CRVLc/OeU4j6L05gesRMpIPPOGqGAzU6XcjDN8GQcVwRjM4s
8GF0rGxx85lN7jDSHDCzpz6uwYeYovsE+cA+TjbP7wsc6erF/4qzgJWWwrwFqHXRnLNtpV62bcSt
oFsuQLeWo5Cb1mBsw811dUQxPvkqVj+5zYZG1w6zcIZTleNraAmQL71CSNUQrHWZd/R45C3T8O06
mdC0SAZeGtdtnfHdLOHpciT9UhcYiapiR/FmYtzOfQMOEQouKW1j1KgSAErRgOZqA/zx+WJTsrvU
9pk8MdEKflSG85H9u92+VKd14aD24HZM6q+eYnUr65GuRKeX1KiMh9ZqsRk+NevwgoJBMRyJVpim
PaWqb5D4aJczqP6hMK+9YciyjWKYWtm4c1e1VqRfJ0grMwNI0hTsnHVq+TS92A/xHtRbO+XBnywN
4qVKW56DpjSrohpr2mTlpvg+ArtfOEFBwItzyuf/6E73tfXDdKYECGpp+8u4fzRwCUF2nL1SAu9N
Hk0DB70idku8g3N/WOLkGR0B5qRhXwxr3BNGC9VSG+5knlxs+q4m3JMexAr9xwsUxhg7iwrZ5m9q
sl/u3e2MTi7mPOwl3mGvamUe2zBpzp46gB6HbIeZFZ39YplJiiekdzeIe/J5fKDydy9jGqA0tlQk
AhcSZuAa1jZ4dF6DTkqEKil+joz/MvYIU2pHswEsr74rjqD3PvdtGLt16us8L6O+82+HrnToDpMX
3gvNr8Vp4kmmlMKLctykfzIBPt0OMuLxYozyT6fF8W64IjWm4GysQEXigwwY1vgSIvz4Cy++3N3T
ktgi6JhaoHmKiKZ7+9d7ZE3cFUrt/sDZNw5qoIoZhieaynpyJn2LIN+PQ8Xkr43pS5oj7f/0xKDS
tJ/2Z5HphNKw68OrL78mm//e+Y2JgVKe0i2TWQxLp6Fb48qZCMBTpi0TZ+Uvy5Un6RWCi20jFSS0
IKJvLVCVnXGDbrlL9O6IsSXzyKk+jRVUtDKXnlyP4G+lkHbsT4y+d4VF00UYuXRbNm233tCQYkPW
q9Q+C5WwjvC8Pcd/+DL6KjxX4MNjen2l+nMqnSxFW63/RrHWAfAujukLdd1iGenve3ibmpdsrFnf
sPFTu60FQ3Oho1qeFVNLGMn98sDJP3J/L9hFfKxZwhxF3DWiHXVxaOm8UdgnGIyZOzBB4f8k0/7k
FM1ZXg604c5WM7y7wiSgG8wZiJ/14qJDuh8NjuFUpjXA4FSWXr2IdAnNsiU+AsAd+/1pkK6SKF5m
kXIEzu0h3os6QVaBETgeaedfj2F/BX3s+VIyV1/AJNcaz+IilarUiuyqXkpJHS7D53nUNSp/tKVd
HHw8Ovka+Jmz67gq17KCLfQoP8JaRJY7YO6WBFCsf6xc1pcxHhp14i+PTbJCO58FS06326sYkZfi
z6xp9MnTckg2h4azneYoI9KZtUqh2W68xiOPghxFKMd2QIrGzqPKn9nVm47AqV+XZApBzRwj9dhK
N9SeLu41TSE5E0zZv/2ratcf4ZNEC5Jd1bp3S2k4QQjtJHK+nr2BR0OVTIV56scjCPlyUkU/I36U
XBxabZkh0aeSQaUyxXiFpUQ8cctoX/+6pHbih1t2y5OUSlB0ga+U1Hqr/8LPkUOM4pn+52hS9q1r
e5dxhS12rroMqCqhZy59oH1BJDBsU3Hpo4TLxrpVrfm1fV9uf4TiRcJyTdxI8cpSIXF/HYmUGWkM
O47CEaq6WKhI39gD0DJ7t88GOrwTcU9Ef5inIBsIACBroBG3KFv08wa89nt9cnNXwbnG+NTCMXkC
jkYlg/Ume4um7exiHlvyaHpjKt8jNAKLvZRxzYAmvGsJ/wTO4V4AvZU84x3PxQjgVzbSyWzXqd1D
bq4fg7vtg4wDXTqTI2f50jNHYyfc92f1NYzJI81dB0kP8I9WsGjzp8BDISPIvtN76u1dv0CzA07/
DMOEtNZU3wYojrsCIrdJdTfO5AVMzPigCOR+8QzIKqw4qjTeD7HiYoznbZxg7qnjKC2UonnZdrqD
Ifj0Ka/hKZiL6TaRTcVABPIqnfc+dRLLAxDtfuAd/JujPQoaEtyvaod7/P0OBXtmFWbp3GgDvCV1
Oga7gKyHVAk83dNOTOP/WMgD8Ew6n1VUijchYAGZr8gU3TI6KTzQwBwyBzlN/XJuPGNTfjJWHpT7
luXVP0QmGnfeghp07GCLUi9XNtJsC9PVzX9LgNevf6BfaNQf25+9eN3aXr/blXJ3VZJcCLsfYDDX
IC8MQddo0DfGSCvzf0UsRAQ6IfnjvVzCFZx23FDNp8VWjjFnV/UI6XTQ83gsyHY3Rvx1OI5mUH8/
GohVVhGx8NmogDTTJ8OkADLZm7EPGPeQJk+iRl9Z02VjikJ0A6Uz2LMXuk6Dd6o0tpq22K6WmD7R
qh0moREythVsuJlYeYNC0FKN8SWa6ceB8Y9tKGv9iabXI51A70bIF+jO6dtqk1qiozDBuilSIbaL
QFuqBZo9JobLEeDyfSouK4Y3P8Fmc+i6qyFbrmOOcE1E1KcUGUYq7VF1RRBCXQLJnTwuAzaeU75M
EP2fw51avABG69Uwyx7mkBmA7fyyX+Zv8ewPPAIgzFMa8JdqL15clPfPr5LQ4XwU5GMWZiJ6YIWD
MfZelOnUv4lzH8B7B14Q+CPMomOSZiUmCvVgww7TmZ0E1kButg2U4CsBlQPwj7PyMorZYbNmqCwK
VDsyD076F7tZ2Yv1eFXV2z3cJTjeRQNx2wuvvFCNKr6Lz9tMYy5uBhkFaBJuWQw8EzCi7PGBRFv1
2tChFfr/SMWe1lIPaUSh2DyM/VOQfN2mINboZz1bAPHI0MMJ2t1tZCqO493joQG2dgCCJ2X//E5G
C2PMG0PoCN1Ue9cQcjnVCgyZD/QRw1FsEWNpK6tcRV3/FsgSjDTIsXwN1DVMG0pBkxm1sepo/gwe
EyhP32y7l4zHIrRjwzUxDBk+jyGWRB4IEQcdfcfrWI1embl1FU7Oscst4136Ck/9Dn0HZv9UYp66
CPG5GzeTML8GrtJHO8882WpNRIkzNhBM/PQNLkx3HGpHAnZsWOzfxtaMxB9srHvvWRXCxrGN9J4D
jgVHVBg2JxnYNPFkFyrGqrUF95HUSFJT7GhwPVsKdCMOJTXC9vaD9X0BWUS/VhKzlQWeD+/9yAOd
vZD31Nyt9sAue6JljDP70M+imtliuaSbsbt1ItC/3OjPmFHJB3/0UPSbYHQNsGD2qCOJgPoz7uvp
e3IiOgfdjdaqNYP8QRlF6nmmBWTPZoROO5E47UxdE5Qt8DuZlQ57Ib3TjTlwD3hWjKDuUfceu4/F
Y5RoHFQIxrPUzwunyUqZcKNrHwBiCWjXkGZd6znXl1lvGKEu3wKrt/Bd9e+tRM/wkV/lc1Ym/v1w
Ny8Edp2DWmeFnmd3O4tblwymD4xvlkLOtp3PuAkd+cpITe5az/95049/UE8UzcRTD3HEPqX2w6Xi
m04rq/NvhC6QMkQtbutCadeEiA4bR+g8QWVg2U/fOdDO8cPjXUGjl81DzWaTw9KrcWmBM5gsxfWV
lTDgl+/PfpmImc8gulCP0xkkNl2eIofVV268DdH6NYGUPxOmJwviuoW9Jzf7hMN0WsNfzKOtaL1T
DmJ6krdgjxW3ge/JLN7dOXirR9+5ak+/fkPnSZkKcN2KOD2AgY5+X7mvxUDy4CbSzndLw3gLq8gT
LUrgQjSodfzt615peY4q2IKM2OFk8zHi5svO4s9ZH6SdahV4IHqi35s2qYaGP7P9qyAyBKK4hjLx
KV52j+P6qZAWUY11s3IV59IFm2Wr08y1M3KnPsVKG9cHFsT8QQblzydapXqZgBL7B7q+mnpsxKWv
uXo7QFt0ugMguAnRk0cPlUmG4gU5Yd/u5SC/7AdpDSfgOmMIe4xghKr03HzSqOEDLSzmbL/CayOL
DOodNVsGwhbVFmEAEgxuLt7T0Yd81FbQnmV1k1lImnyQLN2vcMKt9KDUbBGmlOTybxRwaYnxbW9L
dwq4mwCVwW8pD/CWW6StGSVoVc2yCiOBcsnIpznBrj1mTzdDpaz6WAhxtnhZryZAIFTVsrLtRPaS
VO0SLs8UUBZPbhE2/3BpSfwMm1T1tJfprqJvlQiDPJjYSK4uBh+VCzeTGW8lOPSfrKT+OGrjQyja
3WXsJeIthT5CP84eZgZq0fUEg+Zi6ZjPwU0CA/su05utKotYp27rFhGOt+hHI+AXoRoBxD/57mvu
vfCF2uDPMiJdtCs0LfNXPElYqeBxIYtaZGIDPygHjH81ihN3A05cQLzXisiu8dTaQzhl+jfBNpZd
aErbAixyD0eG6mch3P5O9I/CjGxUik3EM5EJ6bYW+bSLVCOIGy5GPCIut/kvX63pcOiOKVYuNVHs
969Tdc29pjN7yuShm5xATbv/gMj/35hO28LiRBICwbIDxfwE5X8IFx+WeT7BgHDhpcDL+gCxGphu
Cy/dNkJeDRQ1GY0CUCvlQPX7TUzuwB5Im2DR4PNWwfYVASKiBwbcH9QFCAaU9K37b5I+9AfiD8w6
aVMe2VzN5bGqZ5V6O5VzQqtlDTdHLSxBtUsBmHI1l4X89ceFMmUCu73XGXzH8ssZq9HKrlWuepA8
9wZy+LcrDVdHnccGsZkizEw7wNZXAjBHHuVGc8MctUzS3p/4oS0vhyDNuV8hA34hSkuoa/erSchI
PEwK/PQnU00vHVCw89j0wcpgwiBF55YAcdxhCO9z1l1EX0BKyvDZasafh3HLqNVWRvl2Jc692ARX
iBfeBkvDr9aXWrkOEX4RVPbFXbDlHFKV1ndaJ/GKFTJ2fN2nws5dv+S/ZCeJ8u5HZMJsiDXW+Q1S
XoD7VE94mAlV0A9IPlmdYd9ibkrGkmTtlnt2HXWl/Eb2Rklipe3kX8e4bvtR85EJeKmf5XqV64Z2
3SgCpFmj0H3sSYHFOec94l3xuMyUCqxbDXgya+c+GgL40FlVIRpBEZq0XSCrYMVtJhco1ugCgr50
IwJF5ZZD1mpazsBGmypxEhS+g8pqUyN+p85RmwX+sTWkh5b3vBhUjOBWbhi0g2ga1jdVcXztvldT
RCSteVTGvajn+rd+NuTKg/ctKSbpnU4e2Ub/rDjjOJU5Po22oQezvM4guMmCrjrknE+G0Wf4TTfX
o2FKgD/sX5Asq/nyfNNOcylp9VoGsspMR3V4yJK/EKnOEMJRcC3fwgaUlkYgzyGzcCp5MyBNtECh
k9N+H6BhPLeS+mx1vWoKUoX3FWpjMRFRSn/qH7VbCUlz/R8zNONvVM509IIXxhmG8E6k6tuSvMpP
UncGAottcofNTS3WNO+xB9LYxhqAeyhxMUlmJG3/vB0z1chl0a+cl/QSpJTG+ekY9shcN9w7xaa3
wvOleBuUrnZpU9g93q/cs9Xiaa+NjB8ed6AFqKFE6CmjVi2zlWXeX0onEhqQNZ1BzwPEkSx0/ynN
dELBxFKKg3iV+sCvfZDs4A0IGTjd6mnI0wm7jXmpCqaTmzG7gzGCjYP21YlJqv6SKOW83UxdEm9O
boZF5U9YPzO6Jniyq8vFiWfwAdv65BEzUsJemX5l0ZkOQN+ywCbe66DiglI6YxfySNS6rQa+4Zyd
GGQ6LNXu2jgWLyF2/20USYi4o3/a7OO1ARjRzgqVxaPd+hFVDS1Zw+menNsUMuoa61KzqIRrAHjV
+yD36yTpVFTxxiROFTnDbkepUIjq2WPPEuEX7BDfi1wz4DzrG6qes3nWeIH5nacDv0Vis5M0ZtML
vzyuJOwy2ImiKuJ+yfXbxHYKiycb+oHNjlxukRc1hS11ZRFdt3q/WnUkoqPrxU1/51b91nemZXXd
VgEvRR/G+Ec8aUTCLPZuXCXBlu1O+rknVXOiXWFk059ZXpzz/CSwFZZiWkQGOX3QVyHex5lFNrFT
5ta40Og05AECpUH0RzVjxIjE4tVSZw/YxfhGUzi3+5JUtai5oAgJwSW1dciWBc5pMd+6OofDN0Nq
gKRh5u1jmBaBi/JwNbiDTwZieAHf1bZ4h4zw5okzOAhy1DfRmMCTSNOUqSn2bfG1s/81F7xyOXk3
ODsdFlCVg2kOpcRoy4cf4AO+c+0jizLm9G84jRyhmiOpcRlW2R3R/8eGnNCkd0PXv1ES+9Tq/D8Z
+IETmdH7eqINri3mxML4G3LnSsJPtD+O912f6tK0ahdW3uaVk+//3EdIw7B3FPSfOWDvFxNR21to
yn6fkCH2GsPPeISvWYZHtmbARPVYmpac1OZb0IwB+lq2ilEh+VrOu/1IkccB/u1OzHSY4Wh2Qhk+
Dio6Mk6+qTwV+UaVRc/BFt3k4ELBwiNcZ7BVOVK7GeEhvj3P7X/+sQn0U2BAS2Fv2tG5xrETSluQ
trHNOY14rTHltMt8geORj/2LxG7BFeKQJ++JzePxkBmywgyKPMSHLYhqqUfXLKOeVa7K0FfxZUjK
MYVtDetBQtDy8GZtWcDZwH+wp8/yTh2WBPm1k/9vFq8tNJoFR37LLwxtuc5bjc0dyyTUDaIokFBR
YpbdZi3jQYtFmbTNyGMBUhwPTpq1VKAfeY7ofT1rnCYKHrS1OjIj0JVgxhekK2S8liDy4ntTPPDu
Ct55DK5a0qjnR0I7tclQ/hSOcGa371ebhgV609/DhHt9BhXaIReWnsHxa21Lxl1OKxFybacQVlZQ
LfQEw+nvzl6F7n2sQk3YhATs+OBr0LyRoAQXlkoPBhW9lt06tXWC0T11oo7YrwGspcftKAl1bMYN
8af3dzEf9587R+NxWPikAxO+1AmanfN5qRguLGYtnuy5DR6GHFrTzBnc5zziF78QVt1DXJ7qWw/X
BKssT2MxAoZQELZIR3XrmqFNRmOGaEQWaykbs2PdLc2kP0Q1IBjWCUZj3k2gGW0PwdthgqESUJCF
yemhz5dS5IO+IQdQPd8feS3Ye0tY+4WxTqdKL/55tMljdUHYSlrRRXBqx6DPmjvvqYTybpLEVnin
CiykbwAiygpLAiVYh5IP+JI4kgqthUF2TMosxdCSX3cssCxAec39H9WcCW9bSjCdb/gSmfgNr1Xh
nApHMSRVtKORtYh4E+lF5X/zUI9pUP+/hkPYRhKWCOFhuDY9CtyihLr+4dI0Nrr0vef+OSe1MqOh
JajVjUBlAkN6HYxMSLfs1H3z0q7YPKG5IrSj3lNpOK80FLBIlradM5U+p9SaizjJ5lNEPryQ6vEl
OuY+Ru5ftAaGtX0QtAEc7touQlbRew8EZ8Dp4Izv8BWLlR7D94rQSNC4iSLpzTl/QPw2Deuuw+ij
cxEYiwQP5ZKXzbxBhuu0xKGqwn5pFoE/WD3SIUFitFEe2I6UFtJKzXYUr58N0a+D0ZV+cHPBtBqr
eOdgfU2RtXJJ2ZRxHW2aNYvcjK4BahB4nWCW2SLYXGszHZiGqAwatD/ITINJrUBX8UOblLVSzs5B
41tKQxsilqEf8XnBxkQ4ffkSgb5Z6GXxU3KuHBIOKYMOcsKY2Hj5e0Sa8iyJmSu75Y04Ie5EuSAK
lHsWX8ZOW6IDmOt5QbM4z8JDjAbpw14S4KdaE9CogxxnCHx491LwrevzVArpLsHBzemYYqxlqCGi
zAFreWekBmCLnGpYpqGv5TGT2tznnMdC/s51gIsOtIrTwfPSjUfhr8Pr7FMGZTcdbdtsOz6CmvJS
ibA7zE3UADyczzXe7GWcya1BFUJz/4HO30mPIUA1WULqF+KrIdS/IknTQa8m+a3Y5NKW1QVxpupf
cqtdRbLSn9psE+TOBfrBzTYD0SCdmVUHK1SRwXbbiZfwgYgoIHAqSUBmuDuzG84ENTP40zPxTNbf
Xs3qRxjJdKgr+GFBWERli1/cpajx+9QepVV6/bacONx3HklV/D1q8fxVpo2bone5O7wr92WqVxxP
jo9WpfgGBgBdAKBQwMj2RSMENdOXDpvPmFxxm0xY8TzAJ5zhitsA0STaRU1CbM5pMDe20u8Jzkdw
DTCQgKWekTFLS9izTIGHInn4iiDHFaC9p4pMdmQfQgxCXjxYDntOe8ttdDUTaTDk+dJt/lIB///J
/yVtfdCD6Bax4sgAN8oeCFEJQAQLCsO4dsxc95tNYdC33sjQFtAmLvt+npmgq6A5e2oF3VUfLfyS
qE6LRG23X4OVD3pUTQv/bHyTyG7ArPKKeSMYWqaGnuRMXCgmzpD6H9z2JMRzqVoXgoVcD+vR+P/S
Vp0i7iXxU93YFb89UWt+6F7dhBnorRWCC3vUeunNHgloqF47o5aCStwi+hEy9B0+RiF55Cyy91f5
Qln+I2MYuYzr2rD8KHv51YN5v5eLnhNf7c40vu5ycuahGrwocxE6NrnXIalB3fdk17tPJjzOfY/E
pSEHMP2EuuhC+QIoDI3mTwDj+OingU+v2OnXLaE4lR3zheMwYhg5DMtOhxXxO040Mv2kjtJZBZg1
vp+33qZeurojZyE0dMSSDaDKk2ebOMFTXdLREHalAAkbHYEf99dwgbM/UgRyt76+d0yBqk75xOwC
uB9cpHAFDQXQ5XRSwTYzPqRstWWp/WJS7qVZCSJ/tOMWi9OGcFJv3eRjuFxTtmeIGcNJI/1jVWRl
oGzIpa02eemvyj0Pon3xKDzUa80YbPFK4Oyai8mX33JSWGZM0EcY8feHeBILavy3S6v/UepoMAvZ
ASR3hN1hVKqZL24o7JRMR+mX6S4QbTjvDODAn6J66Z5YMbjSlx4pO0nd0qVMKrd2bENN8bLaT7sj
zMLXp0EiBFlDgCYqbV5xk5AfrPM09+ufNJ2jMBNn3SkQOMqgZACgfIQbVdWJiM/dHcJtUVhaqfYg
s+oVdaS51nIrlObzm27W2Y4HyInVlrCXgUjBA9BAF1mqK6AuKHYr7MLVxyGF2lGVcNh71Mx4tPjq
Xesz3Px3SNhAPOHswaxWH9DJYxAzlp7QyDC5OQTKTEcbswhRONT/vIxjoPnWOUuxRVtBb2ZZ+ZKW
WU+6ygicdp03WtYAsG1HuvI3zWJUA722OfAZNB8U9uu/hBM7EK6/JBLXhAsBeH253ecQbLO7NGhd
p+ywOPsl4hIDN51Kxd6QKZt1AZwX4lLlBp60U7sxXNtPlfzq+br2ZbWQPYT3Q8PfrCT7fTKi0U+S
pV4jkEIEFmpkt2Cfl4Jo2qPPz/IF22nxsWM5e7xWaICZ16b77zOx2pSIKRWyxoA+9DpDxskh68J8
xrqzqid3n/OhQYsT0BlDthpQnumVEUxz7Neen+k0bMYnTRXz5N4RGCBceF24bZMT6EsqcWDkWWgO
f+n5m2g77xG2+VmIBOSkcUoQKwYLnjn56ngWxVtLPSp5B/ZzOkxxtrpE5mZakBEpHXDStmLL2JAF
epUcFNesk5fh1WadFZZRH0bL8zzKUlXSCVag/VilKIsnzvYAWH71r7uSR9HrKoxxE5FeJ7nthzPf
kUOvEuJtAYOqYtsfSLyQMbx0LYsRY3PVTRfGeE9ZvdEwZAxveFGCGGaXPMGBRZpaN6sx3TOq5y5S
OupVb/OyMki+Ijztqfm84pPYonRvzbSDfcxwcG8xrs5uBWylDJwsiZypH6s5UG5OU8g+kGlo6gdm
uLcJzEtllHt8Jj6G4j9T5epE+8OglYnY4AEC5YL3an8kUKvuNJjcd4TftNx38AX00CajFYmoRfyF
xjrxYN7Os33a86oyzeDsu3vu+ckP8dB0mz0UeVXnZugyqr7B1bxNZyLwDnz4QP/ESDzApnfesbQ8
pVBi1KMSiYO5KHrFrJuasHtLXzD2oX/inLomVb7Py1uyBik+dtX6GkZ9PvFHrwIYVH0t0tc6jVM3
ZL2QUiuiHkWRIuug2N5P8hc3Dj+6DS54gp4XvsjbP+4atskd9Wb6sKMaTrGN1KgtHZKy/BGRnJyM
dTamPFjMkk2e3vXeJUjCJmrlxoKDUl0q2aMEYHfwFJbFishGpB0KcwEgNEwAB/Si9BMfBA3jZCDv
iAmtEBBP603tUwZ9W28W1QX4cC4XNedyhFJ4OSp9wufGv+Lsq11mJsXQM5Q99BYl8qrvwrWJcbhU
WPnJdIylV17XOO3L3yhHdOG5HHIcrNnZO3A38/MSsGebT0vNQFhkG7B4Ka04AP0hFSLYbz92tChW
cIRFi9tKYTmoTRwrM0higlaAQMu1hi7ftBBHToBL6Q1RhFNd/qFZ34PDaQe1llQulmPHf8TJJYQ6
jn3SuVMrxIqSD4A1nU/ngxtPP+thQhRShAEE9eqyFMlUm24muJiVECSJajay0J79wh6vaNs4CcEE
yMRS8JTtkbeuUd2+58kHFAZlshXjJGg87o27I/4kuvBBzquvgvySqEBuKB4C8OirO/sUioJf1IHl
RxhnQUxuzSDYCabyzN4jZDj5wK5ktZT1HMyMd/vaOa6JJgMK0Glh2zczRglrds9mK/FO1VgSp9Ka
pcw+IHEsDzFF8iRcRzkTCBJaSWKuwBGVqksqEFr8AXrV2cksS9M31eoGvN9FUkTfoo64liTN8GCc
OGbSiMfKVB1CZB8aDxAOwhTh7na3cLp76efz9skMrIq6BrAYFRIAqSZ6z7ZBB+jJQ5v/kKHhf57i
MGBBmb+0angdaIKejFn0Mf5zD6S5LxkGOqgSXPapV59Dv/ExzuorVlHmJERf76jSD+Fii7U3Qcd4
CBWhyQrENo2H1dqItoEniGkfcIqW6BTuvn7gTMR1h8oqiQ9Xl7ckDvlxBVUObbps9gGLPTgKWYUx
BjRjRq4ukqkf38GvuJRYLMsN5SIX3uzwL+3DSNwEG6PMq9iwltHG4/sG3yvVHGlpvIVl7Q1OIea8
WBp6QKGVlsw4mRokgZOOqCmfZNBje/eZlygsHb0RcJcGoY7PC9pWq1AgwfTEyF5HMN8L/4y6jUhL
2w+moIr74wZTSbLl8zpj/IycL3w0wQvov5JMDuxG/6dMYsOeSxa8Xac8e9QCuNo1yRnrV3oq0mxu
iVbl4PTlQvcgJ4qKpQUgqAI7J3mp5yIvCa9kk+q9erWtjAIBEVdU6/A0F4dX4XeSZ3V+MRb5beMf
gcvF+Mr6Z/VkrMcRPT4ZH2qmTolYTCKPt3uEgD9KxxhJR4atePkTB8eqKregZgi8batk0/aTnekB
2ZHC5JFPgmS7CyM1qoPmJTjJsdROCU0eMpLnWwcgQomE3aF9iH3N/5HxUe3o6KN28orMBVBXRIVp
JeZg31jl0n934U84OQCGh0Ly2wu3Hda6cHRUDoPdYwNVWeQ9RVkbErkw1KdVkzP8qQMwXWYbyt+F
oVOE6TPWvCv/ZAAnvYDQ11r/+4GxpDefxI9fhc2+xB40fNxEfdM+MW4ZsN702K4aW7Lr2mApDnsh
nGuvSARa1UFsvxhg2cRT2tw/9wd/uX/VBrTwA74fRSyBhAXZeKiuGt3XLRHBit5PsobLwMCwW2kg
5+bxLigsi0dXKmRqptaQk68F2Scr9ymhLOot8a0xJstGp+yCLKy3B2ASz/205u222WjC4M2+9+0/
YKpI+4QuGiyYDxI7ZZCjIyOBP0SOT9PqePZLURQdNDpA9zr594bnFq96ES2TzHjTct0esDHB6yEg
TUH/F0/Mf8onbttOlEQiVxTPrLQqMTXrNA27Av+cthIUAKztQbHUnA4iWrXX5WrIOOHhjH2eNa+u
yWzwwtQtSU9Rfi1q9jz7s4biRXI/KGl9+Ju++X/qQa26eIaFQXWPfok94O4eMoV5x2JPER0oYVNg
ShAdoHCXf9W2ZKZxwLL8EG3Gwc9QutA4JlatQwZbBpYtCTSvoKwM7KKk4XqTvUOH1X85ZNN788CM
108JJ5/K079QtCmWk/qLkLjRKO1Fo1gVgslRuxGf2P5aei7Mb+TpI3/Xm6CKE2s3w8YiHjbBQFJV
dQFiniANlqW6ZT7GVakR767Nt1wBpZuG90HlT17i1q9IeK78AFmZQJPPm5I8kylb0NZP6BAlzwxU
TVvxBSaumxiZ7vrlxN9Vv6WT2DreW7j0n5MQOp1DbIU2M4shuAoYfoaYpwmwiige3P70La46jPAW
KgXTRF5t2s+oCCBhMgGK4UQdowqsbFYYpTF1P3HFcvE30HxrPwSZlEQdySnD/ew3bycN2ec4PqJE
U5nTsjZ26bweY+wBLRlr/gTOECTjx5lnZJU82Ur/FvA1EoD3zOB8r982KttQXjyT8N/6yfZSAkC9
6icvmq910LTnecTG82/40JitEBIZwm4Wc+lTu/SQOSfqFp2wmFktj7EjWklQMJM8j4WsLU1MSPo6
as4Pcwj9O1VtmA8/aIWyYmQdrd+biTcinST0AxcmVVM/151QZQWKhAXJ4zMFoXGabtZat4GO4HHt
yIOZyWorYJ+2lGY7/N3A7wGpTifww8zPk48eyXVf2UclJLVzI0TDkPWCtc8NgYVm17d1E9Ta0YXT
o17Tu4M/aOSrluGRuGnOjcKbaZ4gnZI/eRz7pVRpI8XZsT0PBMuROC0pNzuaALQ2P+LHRCpQWRz4
v+ggHQ6kSmVJOm/9KpmZu0O7NCKrBYT/zISvLJlOSqt11iXEc60NJ9X4uPdQQ2uPv2/iyYDq4ICA
/ZcVYfe/fcxB9Scx2vUAIU8up+4WkWGaaZ4Ye3yBDVEob4qsbsmJwj+0ZFtBucajEN+0hbqv8+5l
K+hu2sibASRQwMZ+tH3Tpsiyx6gasPOuH0U6L87KqdkiZjwmka3fqM1UMFsMShDbcRPRP+XXspqH
PkBE8r6UZTc4rrsjNSuedm3ItW4k+hFU+tKwzdOSdG8hSAzw78zbX4yGbiimCrBtKbgnG49snCzX
df23n+d+DO+LplNYnrxQFoE20RgXYiH+DGy7geGGU9yFSUGxt8KFJTM7sHJfARTYepMDl8mds4E+
YXixrAwvuj3caHHjzBh1uNgWtntMLh4GqR5uDQlkvGWK5EpUrJTJaBCbwEAQaKIG1bazpxAsghVP
ApwUNiFlJU95SNe+QsXAFIGFm+4DyYVh/By0J1sHkcskrObjJ4twmvDycQcFxHDUhQTYK9c9CrGx
vApzZhP98/8gGtrAStQF/EfcKSoiS/2FKqAR1TNGP22B/PTNzp1jaN+uweRgoUlQ8EhFo681SWK8
go+WTf/ykBw0iUu8jhvrvyGVA57iHaIxIHJVNxvJ39YOzhNFu7GEv8HNUO5QO8nsREEDjrIBQBIm
1j1vV4J+QoNSCRXBev3z4MJtNCaJLDuXLlngNjRQeXpFHMWqLX67TsT0PS9IoeubMSfajIXorrd5
Cb9ONSFY92HzWsThEMluHMhenfJ4ksuLx5iy3lG9cCVsaaZTmGxYRQmGrgC7x5Q2/3n8y0h7KXaZ
GudlPGUPkB0ny3bNBjTmwsm6GRhvTjozNQCorVzbF/1f6eSud83rmTlC2a/5wfS0+sb1jpeEzoyN
510v5JoAO8DIiLtq14wi6qmf2/8qG39SKzZk9ky5qtadRWuy16wripNBtTCVAksgfxB2vTyWv2a6
GV3IQk4LBRuBCPR+WcR/JqrPYJFWo+HfUZUV5LXuLN3fWSRHhqjTUAVEddkptbzlfe5IeIHsw3P2
ORNEB4aKAxwwV2u8D8ha+1aeVxZV8qj5K/a4WAk1Kta/dCZCqoEE/vGZYDv8HbqDhuz2hZ+e+G/r
sKoWBtOsvoOaUMDLOj1W4tSLQ8BwdbPIvJmXI/EushJYRC8IW8iBpze0Ae+hrqIi7SsY6Zky7rSS
nxhDAsaAx9I46sasB9R8AEX1E7UzpFUsXC4vQ4Oi0Kd9j4Cqnig2ejFyzQcKhHisEzgDuF1iT1fm
HtRXHGBglF81qRY0FuWWRyc/dILFKD0aKQj8R7W25Q3qPfDD1LqJODUakhZXY7f7D+SLVK+Ky15W
ihG/de/1hPcA1hxQUQKl6pTk/daDsRCQ9jsaVws/6UXtfmDjdYX23fEEH8AFMvdUvKZvrx8rVB7n
+4WZCQUejDWU0juN7z++SR1+pFkpjrNVw0HtF8I1noDBgjUFu000xh5yzgndrsjHj1h8NO7yJNqr
TcH5H2PnMZAGKG7MlbeRBaM2V2SV3oqxudm5FmlXW21WowEiXMj0cn7SIwtgcPXa1CS5UbBRza8s
mQZ5ukcExi65ETQ9NDNpbDy+CLutnmAUpdQ4MQPNn+AjLMUqecXKjo3w+f/61lsiPzXYEZV3sxZd
9OmU8HSPxYHB3zbQ+SCmWGuYlRxpOoLJbPbWeYngdtHOYoDQ5OQNoFfsp1YWhBDyXIEvyVnkqeiq
DtlZfwhMnX6UONG5aaOA7i6ltPlwKdyTi/DQtiQaozxXYKHWDBb9ndIVx2100A9F00uzpEaJZ5GS
F88DwNrpt2qNAToqFeZ2YMk83jFihQ/hTrxYzj7BA8egGzmCdUwW9cvbaS8OPH78CIX62G75PRwa
shuGHx4iqB2FTdSBSm/lfU8RK5Sek+7+OAuYSJhgLoUIAgEZhGg27A2KegnUr57I2+OhVT35swId
FUK0GUhM/yMO2wmj8x4tZp2+ERf4HNZSvoFHok+QVv5/kykV7qVmN1shoGkh69gQrTjePbBVpiCy
8Jhcn1QQh+U8anS/7w5RZPb/wM4l9fY1JnlrZpz5189NEZcd+XQ9gYOG0RNyU8RO4n0cvnyhClwV
0cQgKKtgUmZOp3W5+gg7UqJoB+G+i4pAbaekE6RPq1P3XfTlAmKKs/NETEjkaUMkLNnbDDxIk2Pv
ibWBTh9lEgo9N5h2wLlZSOGqINg8MOxlIiHAUgIfnWV8VmebASy45TtLSgDRCcu4Z0CXRPSzzGFy
2aSmNvJwkdpnGm5Z0JCTt0AIc0TQtvLxXw+BEGFyAMZuYELWhYly0qUAiFv7Hg7X9zkl3vimEyya
OXbXyJUgNSDXQHpzfvs8HJllNOizxdDpia8lYW1UONYpoaHOlM7C/RRRvyUwm27Nl72xgN7NOlmS
2NTzqN+SviCrtJfOll2t3TyIQYQvviZYBzlfVtbPkRVoFZX1iakxjVs5qT3gHO726iNcfpEmbT4N
O62y2dkgo8CWHbnb2oOtLV0NRDdE1DQB3IM3Dq8S9lHMfGwCZxpRiiDypvwH8grGy0MXtmUd26qQ
7lPnB09BpYaK88fG8T2Tt6nVSAcerIh6+j7UK3FLpqa7I55/XpWJaM0wcPQXPu+KT+1TZARaBsFV
6y/WvSWtnHPh3HAqCKGyAEnwo0u2o1XiJ0vpJgm+tITfDiybLHJyTJeq5J7MVwYz/FwHUWpY8dKU
d0jcwvESklPr464kRNpvAj2GoOvslVSbMWkL49BzerACK6YojO3xuG3Lp6KufTLpyFXuzSoDplVc
aG2qdCdq1uspiTOIdG80PFD57UpN1rCrXq7HRVAsDhx8HJLFs6aKnPowuQiXZyyVtJNI4MpGdx8I
GuCasQ5f+gr/Kn6mma2HdxZSZfnL10+RuUCAPtK2buuD57c6tnic6K2BQuvWrKV0PqylTbMceJNV
3uD9cTI6CRMs8gYIrXDkxWB1M5I+MLJwF3AnK3wIkNQHbzP5vVVgCX21G/AJLrVUlBRqWxIdMw0P
OkkMMDEtHJjwMOZqmtBAr78Bhb8rKO9BQ5j3zqqFaABVdcEsb47l9z28ao5ZnYDfLdsZqBN6uAPL
+RCgqh0i/E6wt4mqp8YCPqC3eY7b2uWtHh2KYE+R+z9+JVYL3a5Sk7G4mlhbhuQ5ewyUtEMdmTs7
XjYAj3rT8mf+o3YZiIUGuXOiI4kfkEjMZ+99LsaphN/BlVdLYZ6DhHdEQTCuysl88sAmgHpO3pb+
XQLzI8tA8qTxILUP18H4HJsYy4j1LYLwt66ENB7OBNxpxGgGOyjnNz9oJs7sR26lvQK9Lqgc/D3J
dptI6d+hF2/0F+UGE8qih1p1xItQs6kmxG/J8l76sWR+8jLlFMK3pz3q195RHfZ/YQKa3BRU8P6Z
vKD7rvdOKL2tpIagvbzGMr+dr+oYOAcycZxnk4en7/RYvEk6lucVO3ve9/qGUQv9c8CcQATVebkp
X2BgtVQZzNBxTuLpBUnahMnZ64Q1HPql+foZ09DhMlwnLLdrXmHqWi2/LBpd84UJwKmWrgMKDbRT
SGKnuPKdD80MrluZ6/2hkZ68dZ5VjflkozToTYsMUUneFcXTnY+4NSV+npzrfBkX02Hf7Oz5JERR
bOHvpuBrkJ6m4wE70mGlpK5ANrjWyAa2TDdn51tA7W1mBXqM0DyYiy13GR2DIvuiH7xf+2s0DraB
FdgRMjqMsWGwYYYA4nix/Dj89IidaEJ2OFwalHZf0T4KDEogJpZTPowr8Kz5GX/dih9y58RKOPFS
dhzRs6VhN1YWaZuY6ACwHiVOP0GaIeVmFDPDk5WPV2mLtlOyXMXlOTek8YUsPy+lFYwZFHYVAutW
dHFTyVbm/HQaywkWRuYEbkZPGH1Hk25DIb3Vh6cz6mhLZaFqADAx56msbiKtfZnjL8QYGQMtlBTB
Lv9M+AaFDE41ypIIdh7lW9/xmerZD/Edk+OAJEl5Z43eePlbIF5hkLLtqs2s0l72C8dfYqBaCPi8
TY1N2vzMkChcMaACdr5E3oAKbRCaa2nPo7NDbw5ka55rlPvyWHnun6uNxr8ZPcLe+TTNLaWSeJkH
nbdisBEN/qpTPUTY/Vqkcfekft28Nhmrfs/b7Ysij0nESYJtzXe/HH74guUUsHmQs1Mjn1Bolp+e
ocO9GFfQV6NOdtvsUyh7cdlec5nI6QLdYJsi6rp+MBzjz0jsOv3hX+fbjuSJIJlpQC2/Cypoq2La
aaItDXooUgYIgE9MBA7PcMbs1+HAyvH2vw1UtyhXjc4rK2FCvplNU1ixmRYakG5t/H7Hdu/S09gh
U/lzUx2Rp79HpLLmmXw782f1sCiJbiawQXZ/JiJcyL5U1b7ViqLDV/5VqA4srIaRkAx7kCDdqVjn
CvdGJ/wy0t8f5f+PX1JUuPo8JMMjmHu9IIuJVUsXDmhOg+ehTD6zG5LaEjRLw+G+q6JIzM22JYoF
jcA8t0BXyHDsIkeaHFLQY+eSWiQuofJKlzbl2+kE4aWLhZ3Z+Y0kWvGDWUk7sfaEsnFJqNvjU0G8
cdrLPnjaOo7bCpbJHvUWF7CAXHw6ML9pqbqYoT/XnWN+5YI9wSI54gUNQUKiGymPueDHOm0/6Qgv
NwQATEVFgnhb3iUHd6TSn/sJPtX9qgH3TetDMoRFFU6xgThWdC/YE3pLSxb4JdiBDQ3BBn9Koj+/
VaEElMuyMJCQ3Ts+t71t3XLKGqfbN/w1NHfE8npvohHSRJDyY3nBVYjxtT1B9+yj/6kGYD4Hu+/X
5mSR+V5bsvOHkfC7R15/vXaLdN8i7tnVYlmN1GNS0o7PrspARkPSwTx363qjxeBoRk3JPyEE5Kdy
trNg8JNvyD8mlgjdNguf7sntKcDDUUfA+7g70x0zn6O9nIz+bzC0uMdhtpJKYVUrsgyl4YOFCg96
lFDM/W6OpN2chJVW6XWTxjfbmiu8rHjVkWNWztc1sfirEkdRoG1lPllJnSANjxsB5op02HaTWSMi
79Z0w6XBZlc9IfqU8WKEjzcVhHrrHGTe7tPL5H8jHSl7fXG0Hmg2qC5FzbOBPvRnTFX9NetsfnIR
HhXBcf50Voy6Ppg2m9EMFDTdF8EJhCle2+PjbHJnB2K61HLctPCth2wWKRTiFan6XQN/nfQOdxcp
84l4iHzqUyHUZVnB9LJ9xQUMLfO8U9OsJJoBv5B7WtUyTuD5hLLAms5CsETwz7TOV6NZot+oCwmb
44qYAUam82sl2bN08zbP1H7SeCYAQF19BjAh82hmD96S3MsC6MMC6QdXN0PlOLhCKYlHiRpLL6I0
olmu2RNG7rJuKjxzDpZ75XHvc9eWh2FjWHszUL9lLjnrjFwrgQXeoTJr7qqll+Ern00/jr5TUmim
laJW/cYCylMVlYjyEIkz+gMqWI/uW4amwF9vvWTi2P/qQy7A3Ucfpmnp9CE0n+iBrhHc3rbP0IQj
+ICA4vCnACgw9oImzD+WZ7ygxTiHFdh8vcKUyLxIDUmwU3b8Eat9G/8hZLKCE7KyZOOU7PeaCSlA
qanN098Qiw2Ijuea5Scpcvzo5kUjaoNxM37GGD35OLaVBMEdfhDesjv7gQbCx4Rki6i6SxMppkY0
vLKyOceWShDc3cbM/Y6e63fM8Yg7crX2MCZM1HQz4/3MIYSCGmwK/0BDomt3XS+tl9UfQnw1myFu
lfyVeoknOxEh2tvUyhvmpXgym0F8FO/TqxafM/WDwexu/FNB9eSOKw4uyXFmPJSbbfWwJigOTwdo
/P6XTD+/0NcXt2I7PaNEHBbYBnENKkbmJpX04FuCJ6lIBAxiBx+ZDXAp82/beCQ7S6dq0VLpO6D1
iQKw1wG81ehGuOne+uB+Iamu4XcSEUBa4uG5z+Vbx9g59ZxRGAEbmpMV+ySDebD0k8DQ/4y/1A44
bVLtltxbDnztEoS+mmnsOhypbfCUAxoVgTefE3Gm8PN2jo1KrNsPSQAVOxevMfFIggH27Jx+G1bq
rYNySe2Kz5h5U4iaxv+I4HiEn6WEalz1gTddyfZuse0GOcZF7YsroqW+xrZgrUJ/c4I83CEG/r53
JlJ0CBTGZ6m0tCUttqyyKQpeVTIdc6+vLZHekHL+Yu9OLK/qmz/14B7g0E8GRyfxkMtQXxbE40Si
sN841wOOAhvE39XYXc4J/yhuciwnJhIj8DiUkmB/4ZwHIXkzRwdwpnBMHPj6ZGG4EKZ0HMAXfRKS
n0AbYsDUGLDymHoXmrbzDYazwwb0YkZaYqTCd7xth0TmKhd0vIT68JzNxZu/I1fgG5HC7rlZO8dD
zgGIPMNmTLpSYjZS5bWk27t53/yGMpJCXAXfgqmyniXoh5vD3dgOr35lzmvpX0YLgVesgfAkdSOQ
AuX/LvRL8YK/ZWT3aUrnG0ht7OsaDyBtxkX3gDqLMXkK3aom5CmOXkBIkTsGd0BxBIbMpdabQk9h
IDgMtuMRzovxueL7D0q+aPVMIHyKFZQraCBkj6gd4W+3PtH3HNjAMzfH1vpJndTEJrDP4tMI3sYv
z0yXm97Y2kw/5070Z+t1x0vK6xnNaEMe/o+Sq2S8Q5Sdsgx37C4SMH79pGG78Ye+VGYniIF2R9T/
S2YbJknCkGoqoiy8RRfhNkLriA+8voopmNOQEFHw9+BYPy+JGa7il8KYb7b/OeLXLYE9da4hCRWV
AVIgphT6oWcqT6uP939HN3z/rR/hg8B4fA/NxFFGGTywBQq2n+qJ4h3mfidajDrsQivIihZtzYV5
BWRu++19PSkR7oO6NzjnYCMx5zBXexyM3fRns+4iJa5xiQQEOrs+TzgzSEDUHjDcagvPegJrceZc
5+RHU4EYTX/iKHehFyRo1votwhvBarIICI47mtU8dRz/lJz9tuviWQEK1TzaFS6G7m6+OpwKJQX/
eR5BqmKsUmfaYRid9bYX6a63hRxH+Zf09gfq82ZDUAvxq6UdP/VcKZLjcq+ZK8ASv37xfKnqwgi2
MBYBvVwHaoQWhdnY6H5fnAZr0fQq7zETuzxFN/hAkZ0SALaO9HSLYn9EZVIwMPwcLnHvoY02MX1R
Jplm73Gfv8XhqzCiUXVrvCcqBO44LoMxA15c9Q30xgqerad9WJR1qLiImIYVgJkA5hb1MDdui6vV
0DCaTD0WnfrGlL5hwx4AM24a+GxGaz03kcaWjozRWeI03ymnovaPqk8vW/CZCUg0JDKrTsqszXHp
ASMQ3a6D/4XLOgUnHpoSMkTV2J7NXFu0fnfZ2pkkS5DFrOu5aUHoLIAabpUlfd9xzW1nNLiMAtNb
tnIHma1uI1fGpcRsWOQnqHVgDtQU+PHG196LPqfGzmvFCjBbp1mh8MIuXk52Odke1Xs7UtqOg2JX
3jD9DrnNX1qBVTTwcxQ5Ku+w7aObF8jQ/u+ZItwLFYDz1P6i80SblYEICc27pkVxrL4AO+Myw/Wm
0U8W1S8qW/EIJLXkk6ZU46BgdLiuQ3hdiWzk1bfHTkGA3Fmf4capms/+Fh00x6O9viIXJJyKuLLw
t+E0S42wT/QdOB9aRPNi8HuuFadgBtGmUWieR45ypMdYr5oSYXHLkP+1Lb1sAv+E2wkr46oKhLDz
lvKG+u6e+cJSQwdSKgZfz2nQe2BLuzuwdqIiHohdEcXXroY84lt6d7LfGK7e5+4Q7VFUjAV70PJr
MH9bFzmZuUOjypYAtzKuNGjYmEzBWQ4fyIy1efthouOUq1lSKUjOPfHTbS9F9BshddkNezhz5nmB
dPI5G1amltVIfb+8WN5dkAenWAzN3X/QxlZ55kEy/9tEe1x1IlM3j9oCOtS7uuN+gYit/Up5kkLg
OkfuQOGyqxq75ucVmgo/QNFGZ8pZiEYD8NROuIkyGXU4KZMR1626AEuApjQtwJHsMM6De9aIQJ/V
zY+h7wg0QFEunG2ahT1n40pTn72/41T0bpFLyDKFqdRYZFKLlGBW0FFWAd9x99P2oojqWEPIFkqc
HNh4k94Ixot61f2ughpZNrL/XAYegbHg2U+FRR23y/v+tNMRpcLMgEtpfDNrHWBKuW9Mo7eYIKsI
PxQp6F446xoCpPU2mRuxBkPVqtjaJAPGN3a1A3XOk25rRiWKbNvm7+LiDWqGvWrUwyypWI+qc9BT
epGJq88h7+XCyfb4tQv9mKJhhMfvm5TAwCtS5tWRPINO6cc7iq2j3mm5nVKeplMxGc1tdCAvlScM
ptkO9Qj/sv9eV/l7Ygb5SwRz+CnO6ygq6rmgP1cTMo5kTkGlmozUNvFE/aOJ6bfPP5RiY/BSiTdh
Lf4leCVFTyuRO5pyt3Rtc3yKNlz7BssHC4EnOilP3oHwVv8G+KU1LK+gWqjOjCFWpTlRG19MbtWD
G88atcijY+71nZMKw/BmJODaS7z7CI6ZPQKU0lpdGLHgizGDD2ok2lHhppVe9Ak4w5nfjnDwXiOZ
dwL6tryCCmIeBkNJfMuRyE6jzWya7wGu048rIo/rbqWgLOvmfD2Dzjqk95I1tGfHv9L007N9HrsG
HHkctzTvDP3tZdOtDim4B2uj0mIs/04UCHrYlQlSSw2eEaHz9SvaBNGM/FmY3DCtcIjltvv8JFWQ
uEDM/QxET/Tl6gSBk21yzthn2K/LE4ydM3hB4AUkwkxxbtQwRRrBiJO/uzImAzYCZtqo4/4sZA29
pwFsJun9NSE2lOrwSB1JrGLN04RbPwGqgXhmzX5FCHsiWKtmPut4nuu4FSquaOX6PIEtoE/wo5rM
SRbLjdNpC3Ckz2WMiVmpjZCA6skJ9APl6pbnAJHYoohYccIa5obC4OamZxyLIx9w1uHZt3TcTxR8
0FvezroL4lDaVw8HSSYOU7T3W6ewFv4bfjBPVIYTa3YgP5fX7mlPMFnZsDKPIa42N/iPZg3aIADx
P9wGSWYuTmJd5tgPup4q/QTqLUVKMBSapVWOjYvitVGugKb8uraT1/6Vl41IzsszKyUhq8Fx4bGR
I0Zfz0PZDi3L+N9TVhce3ZFWZzFHHGtvIZE6VYo0RUgmlK4CnStWF7P2U97sPTTTw5ZsLzcHqwYu
EOVHBf2lwzaMTFzjq2yVY88HIg4BgDS9s4PV6x3E5CfFk2FhPZJeNcNXG9gdgbhCNPze/DL+iu/N
mCdesdUpnA8uKE/No7sJXxkmVT+GFFZG8uK3OezR7kA4oMaGcBcecBtMbNkn3YfpolkuRye+FkTC
M37nO09mxzaz2vceUWZXZ2AQrBmlqtMPwScz0lZd7TRrcprfbh1eVSonigGC+QFyIFuK7i51kLrS
7fnbGU9A/AAu5IY5VW9aRTCZEAf/Y3w3q4JgNYlybabiP0aWcEOKZZbEmljdUNyE4gvGyZS7Ygf8
85x8rV4PBkffyhMgQZH5TSPSr28mXk2q3agKx4BbBQDNvUbtJogQdDUC5swDLJPycVtB4O7XRBcb
qokvIo47pfYaw43cwQi7TKLgo3SWJ0He8YaH+gZS8t5zWRZcBVAaWPZc7iogJmmAHnmND5NiEVsm
qEVx3ojE4fbOMT/H2+2UGQJdINQad0EWPdRijp+Wg/O+gybMrK5MXnXzWUBK9WbkVpBwp5eerfhv
7JhQD/4m84n8bwNwGtAm9i/9C8L8Or6y9C30qxK2hKJn9TUlSHClaif5W8obTwYHpwCWpHRRLiUa
xTapbZHdt74RDOSI7Wr2NtKWyc9EN3g8PnEOAQhZkX1RC1NVoLcJaWokEcRUF8SCi+orFyMIkKDV
eV7ol16xgTnCXhIG0GhFWuugISYHJMWHJAV2jCmFaUO3ZwUBH+wc88Ef7u0IrOcnvekyCLpR6I9i
PYioVcrXOxlKLyFXWLCWQmGe1eh8s8dAmAwtE8RpkCaWXA9p8xDuSYgyV8y3Nas004ji1inxk0Ws
mDt2CcNs6gqyMvG3TPLENbihZ0wNQmQM8A4OlTH/T2+pznqqD54BFzgSg3GLb5rarDTfwntYzWcI
tZmESInesbohs08lqb8jj0X41Wc3NcEjBd+/NznSnRUY3Dt5E1QUp/XLwIJUIwGRkcKPV5CHn2X8
JZOm2aV1k6TVXghSvOrkGf3BrQxFVcPsb64DatRWBJlkQ/GBAKOVsGpscCW7duci4C2oNUR39VA1
ZMlHR8Zzb7ZZns50uN3ACnCaXdBXSSmP7VHSDnYCATFytvw1sYckF396/In/PARN61+6TLEUeQm6
mH23KuEUYozHRZx1CGGSVdlCoFjQfsELUpUDANcAVyafb/otqarVgekvpaXFB92GBd+KyVmVtgyz
JJTNRE6GIO43+YbaMx/+Ux9jY3P1fPyyxWUnPd3ueGxvoh78F/kt4O151cV384Jtgd6HaodJr7C0
31v7b3ys+48epKCIAfF+fsjMIi4HnPcfRXJ51Sm75LePg6BPVvpFWg2yFLzMuacpxDaNCk0yS92L
Y9y5Lnz4IDu3EM6TMSohtPzuGkIgL7tqnAxr3fL9Nx96pWxbYFioVyx7MjazwYpIrAhVGps5vdjc
7aZWRZTmhDLeK7Lo2rFqBD8vwvd0kC80MidM9Zi+5riP41WxPTRYsrvJhWkXNltHeT68eXMkrTly
v3GTnXgQot494o7hm7/LZ29yVk4d+nmtm552dLb9dkjCOhIvvXSJ8R/1dNDTuy1Rsdtwk2/9P+BX
oyaQTMAWVJYjzm/b7iIiBrloPFzi73aTAbmaXCOHgT3Z+VsV2FNLKvpnoDZWoyj/eP2yelJt82x0
aCGao9ujTBxV4wn8F3cdNKQQyBgAAxRQxzZlU6ECCbEWwO1hpcdArcMJEGI5M1JMGRGGESwqBQfo
utJVw+gK857rHMTS84H0tTnaxfY6hBSxI8YAynK23UnmirAJAui8LRmgcDGE6WJKexaKA9VW+6Uo
AeyWqaU5hQIw32EHDfbRr2BiCl/L1fu0SImJmCB5AJZtPcwpG6pTmYDZH4S+YPejHkxiKVE3GR4W
/+yDVzQ6ZT7se/+bkavsW57tjjFFs4LZke49U37vLi1LrRxHxaSEiIDFKH1DVLwB2t/9bZaQOa3G
2iSDLPXX/Nb7TRO1KCelCS8B5Hrj4Fj87GXXxGU7+3nToKzf52fejKlOoyDkOppTC9vMFJd2fu/5
DJV1WBNZz9Lw1DMc1E9U18EAqPxR/tWe9GyxLjGRv0gV2RRcQZxKhsnZsUkungi5UX2n3+HD33mI
3RjG4xaFAMrpXpR6K3L91quZJoKKaKa8uc6FSwKyLY5VEgz2oqxbVMAjwR1qfHr27K3hzgZ9iWBV
w9QHguKZB4uGWSAw4S3803FlIMDESENlLQjuK72NtVdp2Hm+oRjUijLRtFfBKSsQHL6Ty3n+FUv+
8MfIHCS2lIk8vJ9aWHdHVi/FxB+ekGkhiUjSUV+XwZeNrkVt5tvnfRV8z/XFMU3SR7uhZoGcsgww
dYOEJQvNHakLwq6uqguIDuCiKQUc65GDhnPcQeLJmWMy088sz72kUG70/YjiVnHICcB3ALekEVm7
nNLaHwr29MPNQ9wqdBbMfsStl7Us8awhEXoIQgH2Bf3gtA6GNxpJ8B6mzyYCQeStwmJt9GEjcKCD
wEHNjHaVztreY8VbuPPclwghCREj+5njN6qOjTCSi4VHWuJ9jeN3trPDpE58V3Vae9L6j0R/UaPy
85cy7hElFA0mjO25LiQMjj+QEWtoZ2egOWPCeCnOC9KyBuJ2aEOEoght4Q/qs9QDCponm2/mHcI1
VZLv2xfNBJA0++vy7sIWhoPZV6fzbz0ZG4Bvsk8hAMYvpg+L5VgQiVfVfKVN6kJuIrMY0GQqgy2C
XIIerrDPvAu+qZbWss8yYvJgP3TH+zsD4pzn4hT+PnXghrOgqhj3r8356AhcVS/gTuSbpuAuyYH8
+UEEIr1lQBoQdnm4ckTTrNEq8371a7s28mwJoZKoCZBUneCZDD2Y1hWuF8X6tJtIupQoZrsP9WZR
rl1NqsbSSbj+7B95igiESNOcLp4ggBFxPARYrJDRKSKJMauKz86ei4B3ufisIO6WZQn1tmrPaNnI
iV1RMhJTZFb64ByOsguOKz21SVnFsQRQHeZVD8YBqxlq/VRsz42csB6C7VgYWt3m9sJUxvmFaZst
YYoixYUsdUWXT6lYgif6sOZ1QeKYTFT8Ba7dNWOXqD86J/kLIJUl3aTJwf5rhmVuF6l6IqUshIHL
jFhcCWk8xdfmyYYfCMYbnbU8/CErMwL4/a/OfUif+cnxdr1ZMRZu94SNqs0xgW6Ktn07qDSpHu4j
dbQIKQyWXZ3NuUhTegfLDha1/JB0SRIEq0OWkU+iRv/VwUMznDqX42wRII5nOvn5KKKBkKFTk4CR
OOmolnCpWq9IBwoFti/ufoKgD5rIHPGITWLPDpn04pu+wUMvGzmsg4hlgQ9qlrqEs3FuY69zo2ul
RAlQ82sW+ag+Dn2EkvfdRVv9VnLJcHp6/mYlnBwkIBD0sWDQYPC7076vkggRM5mTbttDSyr4SUO3
ChOQSg2WYQUmfiyD9sDTvwyXjE+vOnIXr/4gfd9Gpmx5IjW0LP2+6RtCX2kB4xRfgdChvw2Arg7W
yDScKM6pET2yOMl2V9grfM8KShdLObWHXHgHrxdZSMzZbMEjQK4EIA5AywRNX6MjVZHhdZUIcLV0
ucMilDA+rG+d81RqMHhvWJ/8qimXyAOekZEx88vsqeEdfwdZs+Y3p8U/D6BDbO5wgiuRe/ZCFpRl
w/zpijcKPJlWg2bcNWdAtdCG4m91NOwkcCjxCFEY2R8ZkHaUQyhwZOwcT218gJafS8jbag/DT1Ue
+BMbW9ovxe586BS2vwaMwt4cLNSTm+MoPgT13XmZQEkWPwW/6lQltS8oWbLaH4NgOEjot2pKEZ7A
ZlMVk17/mlgyf8D3xM5Yv5DrBULv/jn1gabTHpBCYoKUiS4hEM8bo84YiluL7+KEvQ6TH9KYR15f
aMPuD8FJMyDiYFeNo/xzFxrM8QZnhPHOdR6gr/f1cOI+lVy8PoWb0Y/MZhvEJo452Uamxtj4uUaD
ESyvTPxTfGYPZUVgNtxnlasHHfV0JI7IjsnnDHTkvz0ZnSU9OELsOkm+95rfOQUe/lxavP60YD/3
mTAKMVc4z/49FWZQ8rZEdzbtgUnTpsO732Vb1Jvd/t83QmZ0Wx1aRO/IubGfsOyE1xHXiIWtT5kP
sDFHXDaPPFZvSdEJ9vruD7GWwKQeGl1G4WRpIEdoOM2nnknMvJkMlBnC6SLqx4bxXt3ZkXivFo90
+HfuyOOHdeqCEFS6Rpyswwtpe9SvUO5TQUBDqLZUQqqmFnV9HpLq608UjqNKekiWf5i623th5B+0
La757YoNiHFbfcgsly0WkHmLLcYdUeX064zPxKK/mpODjoQu99UIGZmAz7tmQyidSOeUgXfw4C8K
aTqRVSodl1UuJ1HHRsR6RFavE8Izixm9ztdLIrat9BGPLAWfUSS77dj2qGvg7TxDiJ7gryGcFIqY
0OPZzsc7TZc0E5g/A/hK/vCLGoo3VuguEbc+AY5m6ExuhOpdZQJsr5pWnjGRnPmCPLN7x6lL3xF1
isxaf40G0NKcioYJdLfjhrngELCfrWvu52v47LJGnw2wo0F1t6LB+7rDETtICCXSo8eKaRjZOV0F
JpJjw2xTBd7p9Nb+lXeFbiX73deCHjQQR7BwHBbpFX/LDNiD8t1kPJm+02Qma39IqTsAykcgR7Wg
TVBwtTW7k2JTIpCyGWxitG5GrV4M4BATyUTHVht3FQcCxe2q61twMb5A89PDkRBmjfMUXHxAPoh6
PcS/ht44DkZanof46Ib/mONDIK0EQl0wp76mgZ4p9/B2x20ytSdBjsnCbdhQmhzLWbDVLSZAnGNf
jQySbq2sY0cYWexw3WULSUyEW4ZC1xAD+MSb1ndsdmms+2j3w14wXEpiKpw0Os0Ms4Szl2lSplJt
X+1p1xZkCbxw7I2YIJsRWxnVJlvKuQroUWVYG+rOViR3Le3R+dr6hkOAOFb3w5rsA5qXS/GS9G7z
eOwObRdZIsFo/ER2TRnkhKjaaNy+68FWthjG6KqMSaYGxkC+7bL+uI+nDfI2Avv+yNPbZwK+DjAD
lin4mFW0ti1KxcO7Z1LEyIuN+Nvol7Yx6fnNPifVWr+Z8SrmfNNP7hfSlSfZ0BRrPI/nEI0XEwY8
yyD9a5SHCzmemSK2pnuBrKDdrlbQCaedtY/b37KHLwcsQ1e1F0R2LdZPjZy9FniFp+qdkclH431v
5c0VHR9uvqnYulxV7sJeDwmSOwTV+yU95a7TgkubJ/kucujmNlCr9p3n5RYHrX+r7+5cSThZvRHH
RfHZWy2/tWVajsNlNHKTnOkyZ5/fziWFxt+bqpn3Uieq7UZcUxN0ZwmWJ/9pMolVajmQPYA2WhNo
zNwK7ZolU6hDgVLrTprOhm9886d4foHG37n09JPjkhPYlN6JY3EloElyQvNeP66QFAfGsaB66vV0
HjFbeYTdFBu7KqwpFZOicVHacbd1NVha7ROPiyA6woermji0sRbERJ5bxNtlkgRVpBR2IOAYRQRO
gws3ec7hrJypP0SrUFkewqxZ+vO+mEfKX0W9qpvLZdWwxcG0lmVVgkIFe28Qjl8fsgDmAtPTFSNi
71X1gGZ5Y+p6+SQxSEi6lyJUIpgtNLkS2UW6CW+4dIdb6QtQa+e5zPlLOpo7w9W0FbqW4UTEbm2m
Xm02j3v5oTYnhPggcsb2AkvX5h5Wys1xa9V7GPO/BFpiHMt0T/I/wOlXh21EsrEjI1t8fNt5UPKi
MO4p8xqlTH0AsGAesBPxpcOCfezpFBKlZDaftPWfmyGz+UgOhhaLSVCEKqyeZpVUMCnRZixXnDI7
dZ059ijtvrzt/m5Uf/suT5Bn/hUech4TzQKgfc87/Ug5Lp9EiCJwyPRPM5Bi2sgKdpruytpAvi0X
yneraWjN0jsBKHAkVGzb9wfB/yqYGNdWfkOVT6YrQxzvqto2/JB/K4rMPSkq+13nwgn397Q3fbd+
1SCJ7dYWVGpXH3MUWmaV+1zQHmo0SKzDc56wNMHevB0Pp0BBnNyZTsUEz+0BBIddTFeQ46eeU8e7
BHtQ11IqvmUgRj42JweYQ3/IHEuma1o+ATWpcW9yNIiTXpZd0OEi7qmxy7OBqjNs65HD47niIzPI
LE9cn5B0CgJRIIOtKQcMmLpGOcMz+y3uSL+BFOkYGg1XHHRbc/dbjsb0mjXxxOrjvh9l6NKa3aTV
OJu0HJyutDbnybPlHcrZ/VO5yhNkkdlqQe4CdLdWgqaLN2tKQ3XvKbv+h0eSE/rGJ5ivAgRDV5Sr
Z9n19JP5DBAuexUYyA3/LG92rpFgVD+fbSCVATsOsMIgacNtg3fxjaEX7P+RAo5YyHFMr683EtkR
T44ezT2kf4AElZCwh2q/ymFdDslB56OH/EVVyZTeLqnOHKicSQam3y1jiiH6MD3JMD9b6//BQUdg
URMYpdkrBb7xw6C84bLq+ZM18y12nmkIo8N6H0Oc59ghKQBJvzSYi53cHAlRkeze8abgVUmsSyvR
YuPZRtu4kr4QV+SnEhFSvAzITdfdRIV+e3vv6jzYvvkeOH6cnds5Z+rPujKVsK+18YmqjaHL4VPQ
eNZBTDVtduvNAjZuxiza414ewpYGSbnkzbBxbdk4JbzLSjIOtAzEHKvqi2kcJtlBH+jvso/m/hOl
4FYEWuxszF8wLC6eLWfqYMO1Vn1xESyLHBDA2AIz47BjCFqoEWk7H5onb5nqSoh+IZQK7iFX2Aje
vO9YM8T+LMKzYgV7i0+Cb9/bypjoK995WTKw1BLygp+hsMIrHzI2ygrd9hEx2jvBQgHYdMns+66d
9C/qceJ1dpfrw93jvIHVXr7DUzta+bDYuzxVZZNA3reOXf8heUlABw8OhGFrvTJK/0goigX+uIva
rIWSSMczgF3lNk6a1AZICto3yfLlX6uMhdYvxSmKjo6BKyhddACUYTxefqZqngK3vDGCUKVVS/VO
5c18qs87qxbp5rwUg4FrDFFbtrUfBvB2J50zb6yM/vbNiMNGTTpZkpXn92KApHJmJ2nXQnf+le4Q
3VQrvTulmSVQeKiSUTed1mrEXoxCz7wMdfmZAzxx3S6KvpNLXMXbsmOlj2L5C+M7yLYBKJhSF7BA
EC7Snrto2ys+He9qIZXdwIaNPkZkQC45IVL8GaOBbHOvy4/z+AxihIAJDvgqdYWTSKSYRgTSC1/o
Be0t49YG6uBqt9yCSG7qeRx7oijAUh67N/amxv9aygZl6w9JdCu+CZu6Y/Ac9abgSQOeC3VI/WKY
yS77j2Lvxqna/lHNw/NToRblj6u0iqg4YjlA496fYNd19OoSyIVa4v+y4IN/bCBH+IPV0GcdBxoL
l6Nwag7aNXnHO4bRVcLoqrAdd1p/uCpB/vK+N18Rtla7C6c+ij2b0XR2en+sZJrVIu4SaB7pDQ+a
aLNdTgyaFNPX2YDhWPLZo/sCW9wEgq+WQCi3neBTCa8PP+BvzegJRx+/+i5chWpL8oiCjYVR3ZNd
g9ZhyO9FuRTIQe38ZBtLOmZqUK1ylVbhSL3nWe2twSRbDu5dMntrnvNq5z2K2sIhe2vl8CSglse1
F8WEhWc+tDFkVD7Y/+fKRZSTYgPyjDbQMn2TlP4bu4vDHKACffAyIp5T6wbWTTK2d2p4JanAheoE
uDFHx4/xYFEcBT9/X4/Xdfzl+I/A9pZ9lajrdv16QP+Np9qi43iPLkPE337qYtGkem5mRbGoS7lq
KVLV/y9vvuLyp/rS6h38e6z100Lcdni7jftm+S8JmCsQ7Tzpd5HjnS6OOZN1qgnOjNC9zIfH6E+D
9kNA0/K+dovNWOiuaWaeIMCJd+V5r7cG4QuHQkm8KvEILVOc2tcpasnWUuNi5Ftbj19jk9kpO0aH
xbT+ccO4nqgUs1C12Y43chZKP3x3cYVFYEFv/YYanzh87c9bhwVQGzm6oVuCwo8Sicu3bmZOPNTQ
x5hB1zBzWC05lEV/0Wijhej8DHavfODN0gMvdd+vpistL2ln1ZQDZS4HD8ue7heu55SSBPGa37S8
bhOWeNAIOBKXCNYLvfS0nuH7ib8T/L9UXdxKhYewy2U0Z2RK169LvJ+Bn6B3kEuhicih1yF1RFEN
vC4ma6HApSmXScjo3wXbugJfL4xFxi448FMIiS4jFYa2vEueTR0o1SRdWqxCnSw/OxFQlUuH5cwV
oIclhcjBiq23RHsZnPO+E6qIQAfj5jgyow6DH3CaMTcC+GToECGaEzktDhnd0bMv4NwRzD1dU3/A
DOWGY59AQ/nDBLqlLJvoM/6U93Z4uljdg2sn2n8xIrhtCiVDcC63aw2CcpTjpkmzl1kQc0Jy2qNL
XaIUWov9e19XpUk57gwMlVJcZcGNnlexu4kK+2GELkjprKa37ai/dLFCMzs62YZpcgLFqON5+1GP
rYGy1h0/nodbLH/fEJHVWLkKPnlGVIVodzghknTCy8QkBI/Uc+5SetWLacy3XkJOaRoYzLmRD7Et
sEyZu/t0p26mtC6O7skthOI5MxSgcOts5yIEBa7ivAlugRSx2xV0863oERSyrsn4quUo74oaaMDq
K5QJo7Q6tcP6LtksKxOVS3xjx+Jufk5V6URCRw2XObMbc0x2pkL56jBYz4tbdQrS9YtZn9ynq2kQ
ddZnzSQxctl89acNhIBs4AMiYS2gWqr/ayOqDraIv+eK50CDj2ka1pjlyMdKscNaUfeNlXoeOAij
SXY/JcFxNeIKelQiNDaCVEC+icX8V5gOKaIbA0Slj/uKEeddZoWOkRcc/S2h6Tt8LjsKbeCD6wz1
2OqpB+VBTlO8CyyvBM5GaVLEx7QGaBiPN9AzTSqK7BEzMZWR0pivV0AMg7es5O3/0QpS/Hp/fBnR
aP0qPlVgK7r1/IAzuKZ7dBNudbdlGpobNUr2qai5vegNy6i+2aR2zMdH4GUMfIxuX6WpzvT9KE7R
Ud4o2C8Go71Ldsv3Kt8d/kLJjn3ltLxi+ZQYh1azFWRAp8tW1/P/YGzaiETIFG7eeRDQjmn75KS7
6nGTj7Th1pmtn7e11djwoIk3Rvhe5UoMotxAwuuf7gY1HtRHC2lEa5QrBaAC+O14GnRbIxlncQfD
I6a18vq6WBOBXS3txRBtqD4gLs2aMsR6zJoPR97GnJ7HTcEMvaZea569C6/JZAUg7vIhtf1BhoGB
bqZNFR06HYTZls4XAwzYmoUfhUTVPlnhg1poiTN5ZPkLzuI9dlzz8I4QdHhHQy/z9/UuGehCC2dz
WDMeDB4S+69vM/iN4U4DdUnj47vUhXXpfdZAl3lN+3Cpubs95JJW78OfxlYuywipr8aSKupv5A64
prisinPT8KdPSIUUb0Y5aA3pPMZU7WTjbqfuYrK10vhIZXSJhnbJ3fRXq+SWni26hpMxZtTgLa8j
OuAGCnR5rekmQVcCn2MhLCoZG5qCkqvdhYCf3ExOLzNDqGCswL3TRsUEK6SL79/uboSBPz9wm+CD
2CnOTvz12PCSukdyI8pjr+rnRsvy2FRq3e6yZC3lHEo9KR7Sq9u8QkuTkrThJuU4YGgyGdVzvQdG
Pf2bSrMfLRZvMKn2jlbFmn//oG7pZYwbk+93pt6y4+Q4rUhzFyTmteddcy4KxkvHUZN32RlEGj1M
o7e5ZLoN3MWhX3M3QRvbnLNdrN0qRdOCUrBTsAVuWX9eNsyUDJ2GM9Fuhc2hFWaxAbPiFb1VEmxj
G+EmTLMp6de1mJZRGTd61BRVGuWaOXpoG0S8HP1R7Yu4j5jag1JOXj0Pf9hEc0/s56Q+MKign6N5
K7b4EiAGWMfpqPL8Gl5Gq3mZVLbwOwlKelgB0uYLESrX/UA2pqxvqJ09hfBTLPNS5l7/KJ/sDHdw
6h5cKlJf4bqtf0/7Fl6O1aUSqUnP3WEUVxY+v+Z8iEHy2brKvHOQ1Yq6yDzIkZBswx0Jt99nF+sc
0lgpH7/MdFE5ZxnWe4P0fwnu1S9mhhQUbB6mDDIKISW01fh/Ymj5OrRmcv7PPp+n+lQ3UkIKi4E6
5bzDXxGgdhLSr7E+oIt7p4E66C2pN94H9h3TNwGCyGH1B+bfMoJXRqABDVa/mPBZPtHwNhRMF4gW
OTirSC20GETZvOgx9Xq1u79vjOLW21TTyrlsamdJKt38y3HXDbbrcy5JFUBkVZUN3sP5qZflhozb
ow1VnYHsjXg0yq0y1J8XtRz1srLSkTfOGWnu626P0/y1D0qizdIasW8Ymeo2Rew43baoDUcHMLxh
XbG4eSnQN6M1uxnrFyBiMv7PGPF26fOuMCmPPfSq+PQbMxkUeN54bQsVhQIfJBNEG9SL3sYfqSuW
KdoY/zTzdYDNdy0jSg/V9AV8usZdFVf1BzgTFEYpnvVtUJcjcc8VHRQrNThNkzXPdlp/UB8Bh6+B
eepL8zrRfLohF2bKNo9gqPyX5O8JdxPzAGk/AVCDbQTnqurK14A/A7SzColYYXCogLbjnhsPpqWZ
gfUqLUHweT4Z4p5YSkXCpuL39iq0aoIlXUrLT3BVUIRiBAi8YOT3sR7X7dxDJqlmdeTAQoFF1QWz
y8qaC7FGMyFHSgySKnFWyOMr/v4xSlJOkD4f7L4DoIpBgQuEsiLwYsbFUmHoEdpu0tA5FVbUutk8
fU9NOlRJyzVowpNQrfdUenJ4cOJ2SGeImjqDoKjddCa+/g8IMK+Dg9lm4OYD23PkqNOOIvQCcszk
U6p37p6ZL6vKWrllsK4x4WEy3Sq8VmgPF3JWuC1HI1ZXm0pV/NqG1zQBBDkLLYoBXpk3vjgRuBAc
vpMf7RzOvAdU0owS5S2h/Ibm4L/wvhNU6u9/DPgpXCWKChWrMgVmSdsGt69+uclQ5KqJXJoirq1r
0ZKZnSpf0CM0lpG7RcBXWXtqEhBVooi1ln2b8iE6iLbiMOmOydru/8LL7mPYBtnWdsJ50gZ+p8Wy
QCz1qRxesTchU7IuiBkS1rEZX1HWgWQ+7YbeleJqkD7C2PELVOTOcjkNjK4Xw5yEy2Tdbq/Coik+
qLW4gmp5Qb7l6phv9IeJ04pWupWr4abwnVinLcwe1P6JKcqYCSN+79ghsS1irt3zsuCTx/xzcbUK
CxVjEZBctxvel5MJkxMJuElT1K1yW0Onm8+7ev255c4VI/0FUuu5IlV3Udc6llhzw6U5hJYB0HJu
A3AFtCDefcOpqiVeAArSgCB+zj/qraK58SYXxB0m3GTv/9dUn23eMvWw9uUMOOXkzM81XmQ+aACb
s/xj+JcLobhzCOZyE4Z2263XPzuZxkf3cxrprVrBFAzSxW7UIKcV0KVFPPVywCAsQafPvIGdKXVc
o0Ri9s8xu9der42Lf2F2kDcuKhyDkDOPaFK10KAilncH0/treYCDy1gjVcYOkhhXzqo89NGh3UYD
YFnF4q2DXjwb58huGENuYnKL+C5iIZs2rXw4IchMBM3z3ikiYN2S9QR8/cyw9f/qxOoCg/g30t7M
wld1UktYKXawZqTHF5yQjGVUhpe68L1AKcOSnC0NVQP+24Pgcb1TEUyFyQsZiQZZycaMcWpChZSh
HLgz8zZOmoya6iSa+oJVPuScx5o8GsEYCtZFf2e0dw3CeJgppJvjc4TseJveIOlOSZZgfDX8przh
1EWM/7Xkg77MBEf5XFm/T1b551VwoM742ZtzNyt0TsTsMEySGRDLnYZG2qBPyqIaiIz5P6YdLhUk
9nbiGSkDR3z4dBcZh2XzEz7bb+JYbfqw7nPzwgkIqAdqiaXkVsDbOpP/cHfHTnpC/i3nnzTb3oRf
9Reey9s4PjSM13bBSc0hMU7yEAe6SKQl8hMLKAqesuJUkU8BAG/zSsZ7SzL314GUoYsPFEt5nBSK
7V+i7yJ1E6Xx0W8evq4yHOhDBqYKn788wobIJaVW+c0duRFgRbcSYM3DJM1fgu0jehxfXlWrESJr
KHUssfuyr+GWMQWflSeTllvr0spR/+lUADkmoAk85y0Lnxy3fDTKSnJvY23jCZ4GaY/O1J3lWX/G
z+K6gr6y29lYqEyuk6tfmUhG4pRUf4W81hj2O1PLgjrC7Cx1kIMdOmILv1qumw2DWH/TUvF4X256
ZfdK8GSrUwAsneDJm9xmWLU7Zp0NgP+aPjNS6a9O5Zwoz4uA1Gq5XU5k2drKKsHpG9Qnj/WVvUvr
2os9b0kHiy05M0VNGjJrC9MJv74oiiSKOZuNUXqGvC/Nq+ybHgHDxLlvab05tWdrWkiBhNJzEubN
+v40rKY+jFIVnPFo5FZQ6DZ0dKNnz4FGGlnm04S2JHUzFYmaiR9WYIdUWQTrvGI5l/BObxvXj68p
0QbZAQjkZcB5UwCMv5wmsvLV9sTM31EDf0sM8Y4zC0Er1uw9AJTb0n25rOSnO+h1LyYIAgVaVrAK
V82ioSpbND4rOK7mPbwVLx3586iQF25kyzOUq1sJG7xRPiTeaZ/9uPrzQ4hdM6wwOUqz0LL7qd6O
j0a/HxLtKEkhzznoUzx1a4ZHf9Yc9OQYkZSknsHmvn/wUzFX2P9amLBidLe/y54lTK9tjxpqaRUh
zvXYtlqIy1fn16vzt2G0v7t+5ho5IaOHPpOdEZ4v66ddN/QgEHmCzeGfZSjU9c1ajYxKBA6XO9v3
FLSZPtZdF1o6VYGC1FuqKaS4Ur+UM82/xRgR1qz1H9q+17yWvOsAzaIwYB51/0xL8bcUYSvgEPcB
WcQpW0MVFovtT7huZgJSjePOyG4fBDsbKokxiz5Fu56seVLGAfETjsADJOf/BDjqsUIQzeoR9mr0
2lTTh9AZT83cTc20VmcE0S/PA4wye3PbNxTKpnrgYJ6xwW6LalndNnF/QYKacxyl9cdBaxayQ5iq
vOYCa/g1/5VMVkrwm/AZGpj40e7kKQi+Vm1XjyhPuvGDll1MV3GPm2vpGSjeNLER7TQGtC+FvUdv
VnAvEkwVvLy/CyjHCLPYEPO305MfgnQYqT8ok8pecvpymoCjXdKyWPTu88+BNojylWExWL6W+pNp
HGwt9fJKZrDX1qg/HcvRtdUs0oW5E+ocekb+BGN2+1I47H6XjrVa+t2UfUl9MNWLDoc40UjkoVW2
hwVyLcbqSaA7amKtGk8znKLDe7FmuhYzhoTcdC4dqS+srNfPXjl47/+8bPHbhHsQO/zJIQZ2QwH9
P4jKRk3S201foYtyWbctUOxMRZxUTMXG1C0BaJ/CVnAXZjPKlfwPloxjrNEF5xHOqr7CSg8768pU
DWT5j58P6X6L7MiVkQ2fvzyjhs2+trYJGXbDpdECNvAmhDInHjSQlA8QEfLgG0458hfXTYktsReC
oXBZXo1k6o0fQg4HfjfozUi/DiOfcOuFT2y7BqHFSctDHVan8wPUaLMmQ5+XUQHMk73qurl7q9YU
9T56Pjk89O66Iz0J39aKT2+OoAfWqQFfdf9Wv9bgwfvB2WLtwU31TBkMStGgn/qqow6PkEw44EmA
4MvIoRNZXosHOnRKfcCRfN3yk4jtQ3WXSfmqgAwxvyTJUN+l3ByNtaLnNaYZ/tRKU/sT+qeNGMTR
hjThybHpzCLx6esrYdcjxoYwkIbtDAD6p51QdK8PjmOX30t6XGcikVramKIezpqFtFfLCxBBrXDq
TzOJ43DWXAuen1Y/dY7gS7y+Jhl2VI2FMWAj1RrZom82QSRcDUxtHrbrvrVeqStkm64q5jK1ifNR
oPU+QU8I6ULLT0IrbcExKaAm2xZL+7yLVx8CcefWH5Yfzmjzm1HDttlsmOhBAOhuJYoS5ajiIQUw
UHz8ODVBYK63Dn5xl0ushFQdmDVXo5/4ggHiBRs9B/IAsoinklSAbXYHdEWLSBewGpQP2mZtF/E5
T6j08q52xbfYzEYxlPMz3NalYna1GqlFJ4LpWohIXA2EPCJ/VPGYLAu22jiqLvW+A2PRO+TRiU6f
b3gyVjD6pxkp9JYmz0Zqnp66C01g1WhLq3b1mFj5Lgc8p0u5yfUu7IwSuqacoKvMNEXkb3DJ7Xj/
tso46axnoJU2ygMJcyoEOqV92ywcZ0bQHQeT+Po1m9+qSGxmGNGkABlfRKSpjgt3OjZ04eYSrqnu
7a8yXH/ipeO0jaa2ebpsVIC6X0JIWJ9iradlJew68FKe0IhqUF32k6WmrmBHpxhHFbcKGhS3HqfP
eLzDbzudxfCtPwxjBSm+hhguTNb+9/FEP9Vf+9VAFecflNbwOBkyulANVKxik/+7gbNj+pZbjhyk
lDnCdYdSeK59bmA2fxshaFmhxJMRFmj+cR8HqD4MIeMWDij8Rj0OFDwRSC9gdchdqP3iBNmckzVz
sRq/TH0jEOxa7U71Erh/gRuusnubDyIThD6fVvFjZj/SX7VNqZ9eqRO9tcdbBDO0k+jpZZ/ptKs3
obj+0lnzdniu+g5cuCyItt64A8dTxl7QFKFnYVbFnC3o3HGPjmlBA0JvlYK7DBFnhJclWJhZzoyS
ZuQYoMGoVpQzMbBj4W5yFH17z1xGu+5FT+vG7XSdRwG/hSep4p+5oPRfyFzTa02TaUEHATvSPPjd
IBJcwP8j7/YB9q98qJE5ZWxRO891kSltIiVW0NEKesnge7pR49k20KE0yQHq6YJCdkJEFTLAfiqU
XDggR2Z90V+8BORgp47qtVc2RJYTe/f41ajs4oDjbNwufK4xoUllDaX6MHfi8gpEtkupadZ6jhwc
iEb4JPLCi6XGomjrSeMiqm7rBre6xcEAbHxaf0veD9dB+x7lK8HsT+ISgi4KbGFwKua3ZfaX/8Ft
HhKzK1wBVqWCgmS56X/5vpSYfldP7OQd9MqK1Htz3SZlVhoxFj2oaxjj7kQtlzch1+Di1vSdIvNr
M6z2bG63KoigXvow6vgRucb48lEDmcH4yfyQ/UOE8v7SAJZMB2bPfW/4ymbjjHF3HP9IMIs8acGs
RDfdaF5Q2fqHezhUZ8MkEBhW9Ye1xyoFb6+mtMT5w9pbPkHDc3hEKLm3GKUWWPbEDS8AnSKxxZ2X
uPFNMljHZOhJnFJ7DOZfV8ehpVAqfwOhHEZB4Qv/K7pu2ZykrhdXPOZT+gO8gAccZzlBFol7yvMf
dLIUF+BBmPgDqo3jOTlO42+2kDSq0G3hGUBc6+9EujzVUqb7c37ueSBDJ2JTcck3f/whdplW4Mum
Bl30uicMibefLe8xf9yb6LItbOrlpeTtn8u90KOkfRgfxammqxG/pbHsE+8ulFO8sEwh3Ug8BouB
oJl4xSpS516j1+qXL9m8uUtLIC2mZll73xqd6yWxNDDz0hEtXW9uYaonNn8y251x0iHUEEjr83g9
Z+Yi0U+moV1Hox+Uda8fQliNUye9gluPlyegRUgAhvqIyLwS+izzjRsjRnYLrNB1u/LLHPKNSaxL
xqarcsUpUx0sUS7mpafpe69jJBT3A3vXqZSPq+5LsO9OkY1HnSzkqyOxa5ELspVs25VSnOoMMHjO
R4/W+xI6DtLdaeSFLp/+xfQwHP3fuIitGhUHRlIpKTKO2oDgfjnoH1e8Y40G8jmo+1pQEW/g7wtf
tn3SevOIzW57bzFK+XIH+00fsprdVAlY4GG+1XcSQroZzb4yGpDsaaLmqPII2ERlcOhP0nXPRlO0
tnFXzvIuVQF+W3CWfnPxTJQTGiS06oALrPJgdO8amC6gQN/km0LhBn+4yESfdoGP96KNTc8IdilF
j2AUccsr67DBIxOM5GGZggdTVLx/zOdJaj0H6XT3UMy6MqpywJK30iL5sIK0LCx1fKErQKSyB7UU
9bz9Hky4aSf+HwXbrIj+EHkATJu+rdVOU6cbttmnWu8+DOxLRguygGQTBEw64+gAluvzxkY82apO
FyX0fvRx1vJmUU3tNQyhUE7KBDu+eGGuCFlqocz1iMtWODr+dyJq5FxlL0C4q45+HCbumJXVYQ5d
qJtU58q/ymoz7FFXYO6sm8MRzQuaIjS08Erz75Sa3WpEgXGZUGtzbKgC3dg5raELa5obteXLkkMX
qC4RzikDpHGTIZ/vtnX5ZStedSNgIenZezVHl3uo7SadKvYq1B90OrevHOBSlB4AuqppL5yTqCOD
YSx5bKVoEoXvL1/f0enEYIvfGYdprQbi3sDE1aFrpzH08csIuScyiEs3H1YgoVTrsNeI0x6gjEA5
ulBPrPvPgVAQJQ57hn4vAs/2Qf7u+npXJiI9HQ5dEISuszgaS9ItYiNuuP7O4GKuLCJagcln2sFl
z3Ycd3vEghDrV86TQa3FY5pjk7V0G+5oljQVOYK8agQuEemTpLblsE6qXiSxReT36BQ7ZvbWwS5d
Qx6Y6aG5y8HDszPdrvx22DqgTXYIwFFj6Fj/83qtNNbbPmZjl0MuP0Kel7VrCytfJ7nyilUXzjrJ
oM+YFXHHzCCM5le6GqS+tyTVp+FyMkLmDAvyny3+Ni3uPAewJxrhQqTmiq3zOm8wtvSs0xYmB5AD
kvC958uGXzl4ablKYvyXnMc6XupA+zxoMbBzyKDyZ5jEhu9GaIQBp7Jc0p0fccm+9NwLVqeqNcB9
00cbTAgGfnDHFYcVwHcZl1HAManXZ/m9E9ra3xPqRV8f4l5RYtPp87ZUQXKFQHyzwi9GlntRZ8Xe
I+z/4SWQ6+MS63blpLGRP2V7jxkuroKgCvoBWY8C5YzPaGH4JMlyzcCTfDxcFAHc9z5UxRwD1wB0
lvK7FWBCWCjc4rIQNRM2RBsb1rhltPGVnRJ25C/PIjRKdfxkO2jMPjep42haU2VKlT+n7aerNqbF
GZo3BYdyFF6Qu2Me6WBjuCMCIOursTk36+QLFFOh/2p4UdIARhb6aoS0ERyyMvo5SeJcc5MtC6bE
gq+OLoYeOVbS8lQQ5w3V5gH4OeJpsUARxeZXen1umK+trCTYzi8oOS1rMnHIRcgYHQYu5wzB3Go2
XJ5gTNGuBo76b7mx919Tey0ibUdZUjVbUW67/W+EFHYKA4u+RkbeJ1wXJqF7zQszjeffBc+2CTnp
HBzq8Oa7WatO/4afGSA1To1ng2E2ygEzwhrP9XW0zML5dLGwxDm9KQPVs5w9tin4dBZ+lKktXyas
/IUSwYDqWwZifSrw+3c21EerMZIn1c71Doekk1HPU3nslBl7ewUjLerYThwLeUaauZsS2i5zrQ5m
IE8rADcloQRpI0UIXlu9vUjbSHF4acquen9eqNspVxXatMilQ+WSIKzoUK0NxxpomFjUdAUVZel1
RMCIG4sIaTRGYBSUO3SehN6fs+7oAxjIRJeq4Pnls94pgGD2n78BHCYLucAXx//rY9sxaDQbxwKE
loBhVFZCneToU9RbmiHtZEI7qhKGlBHTuekphYVBq7u6fv8ppRXvxNr5uc0nylEPGo4fKrH5QxyK
C+U6xc/illOUXu1jK4HIkO/q5djveCOYq22gUcgbHAnqm9roIvHxY0qriyr8G4bnZnD79SqZs3GC
xQR9ZQSBXLITpmV0nUXJ7Pfa1KeCWP1lBbU/o3ZZmk+833eQSFG5XnOkIgfkeGRUYX3LMKmroeyc
W9PeDYZaTKsz2z4frAQiEa1IKWcISOjJGWwTrF7GS92sKsDbfPxwVq+/HNo3cIZy3kpQ80Yfh6Tt
rcdKlxfeed+YbPbLiSv5mB+QwJYP6nfc38o/pfGpQjw1U5jC91LCj2djC1nNtvvYqE/LMTmtcZoE
hSPp0g4joOG54lyTxo5oBXOHgJQPGxsRsrleadiGwXvfu+4A8qLMzEeZ/sWuHPTjlct3CH7xEsNF
6zhSMY0nv1YDD67nnZVBW0qlU8JYQMzCGDmodzRUj+9DRfXqp9dpHf8Mt+E04TRpr25LqXbnHuyv
JpmXJJZ8k7H5+gND4TP16DrH+aN/n9Iu19LrolTSL6EfPkFmipHlGhRrkQQzo4aBIWrn+e9gYaiS
OMQzD7OBJyRifvk3YijTI70FfZ/QlpOWClahm+WJ7Ja4+PIvQWZH6sHuA8blyS2/GZo3+aFZLTzz
unnHzMru7JZ/Q/6OQpIgud8qjK5hLVlUYxKCGbB9svdyx42LgqGUkxj6PVSwhWw700p0wqkX+PYU
70PQ8La3MJfB6cbiAlSYusKR68Yk6uNCM/w8BveaVvE6h0jpHR6l12DTzGSUhH6ADuTRW0YbNipQ
xbTwpcxkG9XlrtkMkvOAhwXIiM5wWptM3YlkUGe08Z5CQCUdq5bXZA5V2VhrdlZQMdE7S8qu5pP+
EQKZN3KzhsMJRTixCGxHiAT4otaq+iSTZd2rcwitH/87o2zuVWvqrvWVlgRRMQsBD8X7KJQaeCHG
sKFj7ujl8GknDQKa6L+JpdDmlbkydS2HE2Vw4f5MTnRHEET4nuvnBheOjzR15oPcQzorbOiuHnru
BdNeZDJw8mcpwt6CUI/OwWYUpxKoSc+DGv0gTmNq9Cw9A5UTyUHmIk9U6M0WHqntSq1MMHUCcVMm
3vBHoFSFqJ/4EnbTUocnG0buv5H9tuqn3/uyXRcs4cufUkcWljPaiBHcJgrTlPuIP6K3FzlSJ89B
jkuYvOCHMzmr6szgFhKbsi/r9/y0epTppivX6qZ/gPXG3foH1CHdAbw5cHxRcmX7SRPv9cqlKJLU
/aq7mrf44a0K1ch+8M5GLqec/I4OFxD94gaf7NkHE2j7CT2fBH2FxE5AFSplIH8bbVSbtDVKE9of
2AN3OuOR51BI1AHds6VR1tiPzTRSL7vnN+0BDvLJWTzu2jRZRDiRQFNVFzCE9Wifc6K1kXVTRvJG
EpW3sDDf67UXQzG6zcLkllL0yScnTN/RgTl/doLSYYMhVSocjjLqXZbjFvDdb+/6PvjqZvD3HUxR
51+Pbmb/WaMExnAiMU0dHkQg77g/Pl/lat83FX/LTbpa9cn+fSS4xFjt4319soL1VHsx4kIkjXWr
OVtmxrpLfps6b0fxbj5giVcYHbs2V5a2aVJoUD8sUZG32xKOeHG/4eMpt9rl1xEXxRDAE2Tb6f0m
Yj8naGD+tvky6qQs5eK03YD1PgoHk4ursNOjZsRGPd9ZHbso8p0LKBNOw6xvxsr4gf3x/za1z4i7
jmaeTNzOTu7xse/VIUcrFdgE8ky26zvceX44T4jrhKxZkPLrUQiEna1SOTq7JjmUEdysHHpa7DCO
P4ByzKnZkQhkxhcaiENq3dyiV4PYpTURkV7uBE3fLtATKaf2RHGksCBm4+2Vw94temmYtpwh6Z1N
DsI9oY6E06KjMi3iy4aAcqtZvzgsJjbP10ypEFlJ19ttXoig6nAMSDqbxK5Z/2g+VJ80HVWU16eK
LVQJsCQMflOdDdz4C7nAgaKUl0wmBpzfADyDePqKNjbxwz9qG7drXJjCJNb6+AH/H4FHnm/dTVm4
DecGfrAgXhte3niKKaqHgK/xdJy8EyDaJItmcUueJfKC5bxrTuJ24IL+CwhVjsgBEVrICixJDOk2
q/UPU5+3OTvOL1VOI/bFTNU2B8Dp/cwqXoZIXpBaA4+VKSS4y3zVPW5n3IYlpnFHJABbpm6Vjlaz
TzxBoajeQNYmAqn4KqkcjbkaUjpa1z2ucvKLoZ/oEBM4BywCusvrORMsZXae2RmfArQp6w0BIRvo
0Dtju+6Yg/6TFQ5eY5InJihLe3lEyPteNty68Korg+uONkUe2u9glSnFwmEGrtHgAiv8gYM1x8LK
+4F6rtR8oQC72w35Zc+63ABr/Bv5ptfOGncHmV8fPa6L6233nBQxSPddLjmv13uz1Vh37d5vcy7v
ZsnijN1mOpjHan+r7D++9q6xw5p/eMPLqtZU9OlOjkKOa2oLVMGNYnSNZAXfRaGqwTNnFzsNeLlk
dyYcMlESdu8PBWBQgdeLhDygtAgrO0unZIhfDllGmhzRZEUt9Ozm6roDPewp/0amqZVixAzzzQUL
laml3LG6s2CA01MHKn4KKUgyNPLARUtff18txmLzQsqDHbhSw9LLZTO0Rv2b4QeNmkSQS3RX4HW6
gAMQiFq5S7hHcMAP3kiC2MXHtvOad/ue9Fj1+JnXUIS+BqYXz9kIEX4V2sPR4uRgOGR75XM87C7f
l6/HO060cauz0T2inENEKQ7NUi9Ui7EoQVbRPyurjYIhuoK6UwqX24qn9jLF6g7gQdZ4Hc/BKWRr
EK3IxNPC8Yh9M/TM3eqFhPzuOl/Ee4gFmEPVyLdRFoTbs2J8f7SVptcVLjM24f9zjHoso1OBOWln
sLali5ppcm6V4O45mJjCrlDuQAW1jEuHOR2vBROzpoI+gqIv0hn8OCz3ozXbarPcFJ9Pw9Bvvvlb
Ylz+ePqZb9p/P2OlnAnM4UbeFus/FKvwRQitcvdlprxS8ydqXJfDGb+avNL6kGeQbvNEYGAgB/yR
ylARC4uhUtStQuVF2Cgyn7jjUACNdaAmuCGljEjXIRolK3EAhimKrdYbNAU9uAeldz+hRpaik5U1
hi0YQP6hi1uKER8sF/J3XU+bN4ZdNwAX3Esa/WuV/XlUJJamhuAkSf5/SLXsGdCvDWNLRwaU/+Ys
7077zONDj1FuhCbnwpNCO5trpwejgq8qs3FzSKrLe1h69bbZP0p4aNFc+BX3wA2VRJBnqVzPpq/1
Xnlx6CbAnvMpxhsNXaMrrvJpHiKkXXFTc+5m4618t8kzpMuj5GeA4OzGVJdwalTQHCmZW7pPBTrh
bhYRcFDbq8O2zbzUZCpXsGHzBSyTCeTUmRwmH5pk1aFJBY3LBVC+/FyD1X0ABUrsH3qLR5BDzaFl
cds2rlHe20zHYa15bXUsqIXheA23MasZaYC6F6DhFsrDqA9+LFAN+3lLMMGPdlpekX11MceO10WR
0dkaWOhgFS9vgPFhVNEu8LYT95RJlxJfUDnL9+kvg2i72hxSskFuwltIzNNqLZ15L9fhX1r/cXeD
HhI5agzXF5Rak5Fktb3V1xDvUY0zFszov/o6YtntJxCQX3ckZjT4DLCS62LPw4Au9CVEyoS3ATAq
9SCDQ02eWCl5gnKdg2BimreCYdoVUAxvExtKa9C3heLEHYjHVRzpNp+rxmYVpQRJd4XozrmGBl1d
OOmzXnwN/8HsTOwpiQ0Has+0/uIrb77hsFRDmS58Wd+TVSx6GtJqrMM6mVQ7g9aiZjBAOJsFzx9u
yMeRXyJR0HJ+LxcqDiJqK8hAeChZv4kyzDNvDEgXaMEY4930BopIrfzT2Tau/H07aiMVZLhZctgz
MRlgSCY6YppqoaC3I0EhkuFQ3S6295OrwkaRsJeARbplmqFYvv9vdLHIG1PobarQLUtPm3YDjoH6
i9Scv7MeLPUjovx314LwTsoDm9/in3Ds547qBwQ9k0YMdtK3vliP5xfdfRKG0LbcpZz/SuKzeltt
MQclX0TFZEb8QuVRvRV2pUMlS7s3lPanXz0lAlyYnL6imxvu0ZIyid75fgU/vfnXk1n+KAVqJ5sy
bYLSCl1t8K9wbmdZJRg7kPc11Az82TV6M+/8VCQYdmVPq3DebNYJwmycigvjMPvdNDyx/IQZ+xm9
bErTIsce1MWY5wnrjLNjE+0DjqCTf6X/HiPdH/GJPVQqGweW7cW7xzE75GkXgleeeADiIAbY7Cmo
VRVPDP7OJ7fVGUKbhSVBtprc1hQqkK9LT/pY3CU5hITVBPuZB14e+VNDWT90DO1WvF+R0B+JkiIo
Sh7DU18l0hJ0STp6w1W6Qs6OOIcP18BoFPuMulm1J07o/QMNe4WvIyD5b5n2pseD2q3C/GNOn4N9
J4Z6hJk8ulJpnqqL3nEMAukMVbBQCbzah7Jf3VM5NikHjcfOQBIvDVbUFmTNiO/hIejfspCQXEEV
E8BHxy2D18OY6T2xIC4UrdAW7L3oo8skEfKpUsxlh8+3LTb93AGrFWTy9WsuPXdw5JM+UCxdRaeL
wSDtQf0tZfh+gi/dg+pAKRkXUg/opZgNO9RBI272F0YYZ9soETGXUQsv1N/+q8WEGduDq2ZfOOH1
FMfG0dRvJ/uGWcYbDL6AdCZlr+PTsO5IeH09FlTVFxml30obtzge5c6eUmQE89SQMcZtcsrSuTZm
ZfVN/GKO3Rk/il0uzR2k3zHuadeglf3kUuzc+7YqYDaFFFb7AXvUY79USB6T1QzipKvgh8SAvwcw
nzJptti+6OMtSSIzNFJeDRjrtEWYhW6TC5Cec5pR5WkAPa946Ua9cxQi7gyqoq53ItUe5mz2jUoL
goQBWYCxXwH3scUWqOmr8sbCXJh23ML5G0k6Jok03nRh6EOSInKZ6Ii79FgSBhBzeTaXzHRUjfxx
WESCsBGIAODE90jTEDYGEstnw/aKUh8YGtDmaM/cKMm4DEg3ehww7j4xjkuk0SVoMx5GaidlbpFQ
embvShFjnH1CWqdEBpqsHBP2rZ6kaD39u/nmY4YYo1IO7mWaRiL2IrIx+gtgb957lfiekqDBx3IW
gX/J1manfdvPHoojweTHK2Xx9xva1YYOZh2zB/GxMDHskqN7WqcRLU4Dts0cWnLV2F8avo5xP5zO
Syg4NrTEiBqiHWvanH1v08G+kW8NoYxSpVp6OZ9HCU3vc3Yl+gHlvrw//0i4DYeGH3F9P1qtpN+1
1eW6oUdgPkpzJkNllECmIOZtBsOahJpH2mbAqRTZGrVsPPjP+hxC5DbR6PHcRrqjt6JjSHhaMXNp
Z8NQuujNY6ZOKliX9lVsoyItz8M0hiw1QLcj3Hw/1tH5VhqDnN7aNpxCr11nJAMRR5OmZmQIQFoi
X5VwLhamC0jFmJQ8nlV/LY/dMfQkBpuYm442G8U5nW2KDum29JeGnkhee/fIe11VZ3D6b8Syj/l/
zaQKX+xOCNoAkgmQ99NYB0APNrvP41mPJ5vCkJAhK5+lgiq+PoKh8tmcCPcgz2tUGJKDTPZNCVbH
4xsyWh8x82bzjUyuS2ZLUI+vjjoxivI3f3Sk8lUiT3dwXeZpNHj1s8dGqq//jCHp2p/t2H1xGefp
XswbbdWSjy0coq+oR+9Ps5XU3EZ83vEYpWO38A8x8yMyQbkwVT/FJbfR4dDwsEBjk2m5mvtAkEBM
X8rdmvjgFqaa1d9opDtBXz6vpH0Bo6DPAlOI72sP+eohosj574yEjql299W58IUsHI6RlOTdSStX
kkVR04ipaRumIJt4MtQcP+r/yaGMwntE4hqS41aFk8910f3OxYP7B1k+Dyh4IvXJ+2o6nfqk64Q+
H6xCbNrP1wInLokFYrNHpxdOvtJaJeRpRuCNun/xyv3jHR1nqPZIQvkr0ioqmeJiJRCZaoSK8+Q+
Ue95j96giB90qzrIz7dsxM9TVCkPecv+lQy5bQXRb5Qj550FEqigowvS8ki9SkNhkTOhgUHtDKw9
b7xNvmJ1+oFj9qJMeAeEa6MXW7cIE8qcpgsW9yCf2bSMPb3dZ3g4EyDTAZXb36rIisy/+NY6LBMV
g95KaZCqj4hSiBSZ9jTVvvaN1SZgBHch2fECHHloasbGMUhXrkwLiE378wZ5nBLUUJ5dDVyXcVWE
bg+wsMU18hUxjogLBSq1B88zFrr4v9FvrrAUnF4WNfFWWdc/ZyfkxetsCnBNkqV/UCe5YV60oIfE
sT1wU+ZQ476kLrb38enEBQ5Qn4RV3w7j22GBgm4ayNE7aZj2dGg77RxgpAouLMtDcQeJuUn9FOmA
mAYABEOJu8K4CV9yIlb7KJVtn3+kg6ctK8/ZaHmhQUPUqkYfup30WNqhwUy5JDG457obgCcs81YL
LJxMXA5SANHBxghiD/9XtHzyFTWVLLtrC9Nj2oIZTIR/sjIZ5DMrTcgXeEktAr5PCvH09pwcrbZf
kI8OinZdGstb2JiqlMaGhFmgmicxeKi6oc4rGpP3G/XFPysEWeezJgTETYfFuc0PSEuNCfl5g8o2
MaDvIXm3U9AdX9yelc19npdGRGIIrFe17iFwi7S55peVdce9P7awoyG66Lu/0DjPbfhEnb3E5cXx
RynBY1sxFKwCJvBwHkRngFXICy0yqEwrspSU41bCvmUI/yKvS0kjsYJSnEiMtsdGcsUQSSOI5KgR
DMRSE8YyoAMit34DZHgWyiHIUtxfMyM6SE4TJ/08OVcdmdfA5nlg7Y0odwg5Dd4VJ6gMfnfe5wYk
FpKcwxxkCtubbMNMql8EDrRSCLLYhDHxVWqLPCv2FwaY64ThEIW/GAf8r7dp2uO/kwfwO2j0EuFR
X59KRbhXmKjFxF9BNbKbVAKjyvsc1+Y2xTodFjmSQL9lJZUtOms/4bVgObWHLDk73DU4jvCyBVVi
IAfPJQOzHrxFJmXSYZQkSkDUJTuXBztPIuUQ82E3+GiGkNReZ7vNdA6X8Gf/T5KGZsULFtPXt5OI
Y81GvH8Zegm2rY+RoDNnqR1WDoq0Y98AexmWavZ0NGfIPIPHxhYuh9wJg7Hft/AX7eL76DayCqhS
BdDTHeJVodft4D+7GE7UBzQIFdr80JZyQACD1asWSUqIdnQ2FsX82Wr/tiWW/Rog79JGyBLqvcyw
7odjq2sO6wn8SIOlU+doF1DTFwyUnOqMEtzuju6MtLFDNA5ftKV6KhrXIVqF6vCffhGCrM2ntHEK
y8qMfqd/BdjlJF95z9hUu7gP9j2XCU9MmRCZdQemsxzteFjD1TXkyafaM8Q1gSl1RjAP2atUJQml
Pa1lJbnBTE0F6V2M2F0FbGzGWw021ZlyjorzVHOFgr0G3d/a8cpHQN5mO3P8P6+2fK/PfJ6ljTdu
vtqTfRuPzCDGRrin6k7WJDHDTEj4OuBdPc+z+f03BMirF1BpIBqhc074PEGtV7xw/EBw87XITBIb
6e6OdeNtZ7ns6t0WFzBQ9tOYcvfEjWaHIuSkoh0YwSS5r+HQciDdO1FKL0SwiUVwQPyiSAGEgcNj
r8oEtXEjzfg7ifJlpwayofq1d+Vh+mDOHqQynTcz7MMxveOf1p5Ri0+mPVatkFeaOXyxZNx/4E6u
kXgKBmIcd8RNMu5qiZenz5ZizJGp1xtSuLZa1NSnhIFvoctMo7ZpE6Vm7KaHacsDDYxijzgPfTxy
+QIy/jnYtKEdN7DVZU8pBMVlA+DXF3L706i/MaY6dX1Oj1JNPdWJ8Mbb8ewLkPtba12//+GWSPUD
qFerA0ok8iAW36idRYlHTuAq02j3qkyLwlzz86heTHv0myXokJNb4boRaaP2LJ7mpyFOMlwA/CvO
ctL0fq4DYPwQJVALAjo7NpZMCmCjgye1zjOKNC0eZj33q6/DmAVO0TRxphClPS3lSecJS4fHTmmF
YyoAoLyVBZWxodNOPXyEmKxToW1WTjmV4hdPah2xUlqZ8puen8tU1nPizttotJXuGJ0B4O100w54
9eORHIkwN8Mo1cyXoQPFxsyCmWdZm6famyxGrq2v6s3mFSHFVm+hHFXsQ857M3tZEzfTRR0Dtf7B
Hx0g8ZDYLVwQWrPrIdfdAe/CedZS7UyIQOOnzhdhZ1QZx1xC8Tgur6XpIw2a6N87jUeEyMf48CFB
UIlTxeQy3x7DKtsqOqQReA3S2HUS181UPSHJ8LXlnbGdaXZaHcRfbO9BAqjcWdlD3ulocM86sbsZ
Cb1Oouu/Ju+Pz4BNcxKETalpLfeZ5R1hfgYKwoL2jhupBsYLhPARkhSvEDxBj8XX0Zb9r/oyM4aX
SoR7BEZZVQok24IT/FDm99X9iK3DFi7LN7SLAjNLK6L7+6/8k83q/zP7Z1TL2CTG4qFRk4mbr+8W
rScKkkWdZ1uiNxQ04uLkYJVUXcXjQDibAkQ/MG0mwWbfRnBMlbQWa40VDqY7TfGI1YYQkT3xbxb/
CLwfok51AwCe1dSD3PmkIOL0hpfehvQAHDDC3u+ySfVZM94N+vcbF6FnILHyGg/t5lm6p2+x2pMH
NGFL4dHjRsG+xzk9cbGoifPT/czgiblONgp9Uof1NtfTVakHg0x40h3GWA1FYWfgIhoJvTDmvn59
NzbuCKpdTWHeUXHTzfbtOBqEcBpll/znfUaKg9T3qoGZhttBogGAZ86LeU8TzcA0ULQnVLrssTFi
w94oziRS6JswmElbeJMjutkHXaliVHIj24vqnBW4hLXC9KamT2PwWKQB6RE4Gpb2YKMrLwlaVfkl
5h5CyH/6ldVJT+scHMwZcbdVuafWqQEXqX8sVKs3gMQdjZloVlOaXwDgnL8u6fnoFayUgfjVaLKc
sxlPKHxT+Xe2tE7pMo1GHRvkPRWez1THXZSRdRAPDqn5cUJAFz0mz3dAVWH1rzWtsRPSBZDM5LsG
On490ulSDxFCMqADfJzpVw2BEnNQIQrfBRuS1SNATRVWmVZjgKprLgliw8leKkECNO7PVIVaaprA
BtDVwFQm7zPudI5TCezgr2Qd/EwnOZGoaKmcuft3KV5NYqvyZ3iGTQa/MAOIbHCiNEPvXvD1fOo9
0l/EtdAMkrlPJ/bl/dJnq4TIZ3xPRwC5gAwm+x8GwgiMlUtsqIxi1X1MXILEst3ZVIV4D1t0LwTB
Ms4P0+RUdO+k+5PX6lurH5Dt5bM3s/s9nC/UIFVu5xtBFiPTDkSGmS9CFFDX91IN+j8ydnVIEgib
OvfySTW2mHrvJUyNhh8nTt9bJ0Z2AkYACicW3nhDIq+00Y3fw4h9m/+d27TlCwqzJ0tEI5ASjKBA
4wsQvjkqrEhmnMzJUxadahZKgi5iWNhsWIHAKueo3a77AY7Kg+bt0z5fe6zuE5nmcpU7beHy4ip4
rqa9JTtRSTsgtU6F55F5F+/B1Muq7sjzXkUxJkGzSgm+uKkcsuK2TncFlaNpJfCRvdhn6pT9DzAX
/OR9kdBDzSVTHYXdlt1hKsBcluEaPY/wdcSjD5fPnKLu4EabfBqW9n2bTkhJdGlgv55oBCw4oP8q
Sy1zTJwu87E1OWLRHDAp/N/eIK98/4LI+6iV24XOraQ00zx+jEkiNburWqYDmTMPKnUF8iLnrpnk
EixHMWEuGTh7tUdeDzF1egRcLjLBKoKqLxfxNOoa7kMSVqcZW5KHr1gZFQgzfHqG6Xe/p5Yv2XRr
xRbwz3W2cThV28AtoqeRyouTwdLHpTPFxjFUfbXOl+wFNGdxXoDx6ma+Blfs1nUZmQ/ljxh2e2Hg
3nowFZYyby6zvhpvpvaQOY6ULla1Y54sH8M3xlHbc+LFAKIGpcgENCS1r4lUZjfLMTXGR3FXgYIZ
I4nV/vCUByQVZ8E4UZIw1cI4eI56//5UIbJMYh3A7u+qh1pHq24YyIOY2iDEIVEPf6Z3m7MtndA7
sgVG9vgNjTtH4WUL79rBF9pkstIH6bhKX7SXKqFd1tLq8XfcYDA/WKMDLDd9EQJTCg8c4ysdaNm3
/HeMnFXAcSF9nIqgC7kMeIrdoHZXBBJtlia+OPLfMGZQ0Ha0igbplvSMJn4Tb/HJ4BU0z2tCrlVD
ToI85+d7DWkZhfS89jxSZifnTErQj1j+3pSSOkdpHBO78BREOEQfqYpVGuUE779yJ5ewt2tOl1mD
dQwrpU6SzpChrjhGwD9m2IPO3pukN3CmvYnfDSKgL8P0C8G+MAGS6nFa3lZrUyWag9e55UxvtJGu
WTemoOmLa93gp29cNn/RFQA3I5nVgXFVe5BrS/t/CPiQSbjgONw6pwF1IaxuVXWSuxMKZou+/lSh
qqneM3RVYp3LBzUV3UAxpEQOmHyHMJ324xWKa6euKU/okbDZ4gxiyntgJt4UK1cTpz2OXGoUu1bX
8dqFO5sh6CxoYpSn4k7CbDlC46rGkHImdXcO52zN+ohBwQWXjNAC7RqQxYu+L3r4/XXv02TIbhzR
5rMHYFYcijYDUCyWPjH/tqyfGkwVTHAwC33Mfv40VFFbii5jC6XGKRcSG7mzStwCEjfBojWy7JS7
zUQKBpKNNoOV1KCcqtMd1IdJ2msYCBo+FqYJMClAxeCQrl02jHAxBhzlXVJvXDh7966iq9wt0qi+
8WCLJJgjn5C3PfOpLyrpourN7tk6mPqEwOIuVTpmbs1eHypyXggK0LFFs2kSx3y0g8I2fxu/pRkD
IuRLwG6AOR+N+zQwg2e59MF9MYgimdrpbDra86HgHBuFDFtRiWJmWvRF9oqzNoTeeydKxKrM4mAY
NNc0z/NvkapfYF4oe2AFdjNKacoCrhkSvgslCWfcGisLNgK/em6oK82z/521/VUgQvH/y0V+e1pf
Zo3XTcL1HR4djedeVj0jtTlJ/+kfm5ajGl+EdG7fjekOXG/ix73oKPmsL4xgplE/XB/hNyi6clVu
x+PMHsxPStB7FmgUTOzRXzHdQJRXsjaurqwIgmeWsYHTuMNZ01DoWV7iXur1fjr7iQbsklM84Izm
etGcOoAYCOdkCJ06bD2BfCXn9WU3w0a/vPEPyeEeGMeahPPnLpJC8lG4Qpj+l5j7T7ErJIWlTuTs
5Te8Cei7n0uB4XBGrecGJWe2zX+XqgeC+03+F7qAtOxpwJh2aDN7O/leyI9u564u2RhMuPcysicX
rpnJ75db09gsreiTDDUuY/FTPUULor8KBseQxAnzcf6b0rPa22/oZjUuMZleuiW4vGfuyKbz1Dcm
FGAG344qoIV4kBSmFJDQNrjsxdjOZNII+EJZEpHLnSoFfFl4aO2HGzj34/dBW7uvX+JWoeQj73ux
A7JSOWtOcZYzSrbfpr8VUYem7QkPB9kc0sPr3vvTNl5jIfts3usxt4eQCLSjmS9h8+HmCCx8gLMr
sDSLhzsQyFKwIC5A66oDceumnmJIgndlbK6lVUQbgUuQ50RVPlVUZa3r8UeOnc4dfQewtecuzhFx
/C1d9R7VsDbhpJJ9VBfgE3wq6BMMbEV2rHEiq8v+KZj9grqqAUCUPy9lGo008soWG28hnx1qH24e
oHmYNjPcCgCqyvYtrS2MLLKZBaIixbUHKHkyvzjEaYMXRcO2PxhMTSDEMB9/P6vrYTlmjs+GwCSg
PAd34p9NTCcVry45IEAs8mJ0Q2Aot0tE3n7cCrX17t/5lij5ECwJ6ddHDeEpxg/bjOP3Fl5gpvxb
/ZJcQd9kFmndbnFo4GDwfURQdnVBwAL8fI3MAKnYfgMiWbyCk6quu2/i8hRKH7EAk+8LmCTyAJ5f
pnbhvn0GU3y2n/UmgkpW5uuVU8YUUaG8Tyv8Sog23WgrgMebXS4uxlT/MbspUmAdJi7AFp8+cJ+Z
ACjO4tOi3QB8vDIyAvJLwJ+PuuLFoN83wvLpKbDXfCIBTvNWGxP3f5Kfj6EJK2O5/ebXbm1p6eXq
bbvO9gBc3I08uNbt8c8/wBb/R8fKvAqls3484sJV/5mQuYTRkZDN2L/MhjDngwEOWFdWa09vd2jH
rceTQKPtCdZg53reLQLvwQ8eXBwvVmVF1vocIfqVS2z+KRF/EQtzXRD/nHG7QsbHJdM737mC+OJx
/pleQ45Ip9/tTLuh7xqdgsvd0OUIEXLOqgvk/Y1pfiUgZ6mVMcYFG7aJqnfApki6VvOdWFBLO5Ay
XCnsLJYt1alubpLrJiZwE+ZNA1tV9oKhHIhtZVV7xSJazQ6GdeWxb+gGh5tHn/CkT5Y5rF0istee
Oc1nfx0pZuUJs4c7c9i6DIuBDEKwuokgxa0/Tc7+molSos2UM+xLpUUBtdx/OXzxNx8gLkyqh5Uu
4nuZxhXS3sA3w999B7UnYYAy26xAyIbnoLylT7SW5R5n7OKzV76sihiJNIJiOchdYGkK0nqiQ95z
+F8zuKYTJ5Owzz1R94EixCNV2nz0p7xBGVCB+IBIFlM2VfwMB10Y+1auqQ6bRF02lO0Uet/CRClO
yJdk3E6KrcI8qTW0wJ7AfnOU/MXIjxjAHT0S/YSr/mKknJgvGAFyuYmsyDgzvaHrgqjHMMOVhcJV
9FYHAUideZ1JLyzvQ9keqWdtwKbWZdGAwkCpSAXChCQVfCT/PNmrvGCS8VEW3NfjdOUDRbp1tduQ
JcPid5NlQVkUbq9KA4DQuvyQODZKR9KhqWs1LsRJysk3gy0eY4ryhO/NT/uoNr+dPS61laTjEuO/
vrpVeaytOL8rDjfMO2lQch9s790sIybyiBxN+anl2kiiPgit8StTQTqAKE2e+b2wqjRmgyIDhzi1
t60Ubt7yXhkIAUycXJm8iR7sBqjWuLgJ4sBInCFAbU80q2m1zrKYINncnK0TCq5kZ1kqc0wgdSnr
w3eFSYVbd8Nab7jEPXZ9GI0bKazVt+Cogjkx21Ed+6tigQ6lF4vP4eHmEoyRLZMzlO8lVlpTc65N
qlMEcggZsirgeNjUo9CoLQiRef+TTuLBMq3rajUQWmJcIn5WvAoiZLd/jsxZp5WxpzOyURMp/NUd
+tPJow9Ucp3ttEJeUMvT4VvJEi56JcZ+vNc1MaRt9+xsvrixvD0EiomREzatngknOg3Igp6y95+B
009EvR/Q1aFef11c6LScXC7l78OJ9gY4z8AONgb93JUlxOqv2N8ac8D3aUMZJgBEIuttVEQn3Gag
stbYi5xwEz/tK8WJ3hKsozZBm3yOyI8Xou2eShc4nMF5KhHgez52l3nm0IvtAy8u1LQWoobgb2Mt
kKlQvsZim+/qziMCG8XtYQQBLT6accuyVLuhcY5P7age+e+AfiuG0b63f6iOHBJ93pBYNllcGAwi
ERd1tpbn4yyO0TQU+Jpq0Ce+O8BgdvRmEOTLs36hqOl15ykFMNeNK15ke/PEYq88gTRpeDskvpeo
LFb001z6oU+SBIaHCnJ8QUflYSFmzbhAqjlQV6RmoMnZoWS9HBCiXg83ZOoc4CSA24U9k/vd3aNj
PX+I9zBEb+NAtVZ0KL1cMzYoJp1JXnk8MuIrdy5vLKilBVzF71KwGNMifXnSoM4nWfxU212CrndN
SNaw0b1NvHxaCVns4DUHvipEes1Q1KfgU7FyvosmG9IOI9caGpC2zX/x8g5QBEvcokgaGTfvEgH9
0X5DBdbF+1itC/jw0SwSlmy/ZZgwYk0q1BxgZ0dpIDYjeIW8+78YLbsm0uvUvS6e57Ua3O5ZruGc
aavrTD1RGfXyZaiiGAd0MWL+Z2uHJbaH2W+D8hM39RTymEHvIgNo8jiWbDcCl9vHfU1UH7P4aAcj
LVzFdqnlaDjt/iraJw/HrZimefpRof2QR3tl1KxJYndOkZo9JgVAcF1EJMkgDSoLKHjY3MPP3wfl
TecytIcW7GACcZt+ExZf18IY2Nazt6TXONhrSv8ncdS9AiDDo9HxUw3IZXCojD7RcY2Vj54i2agt
uz14VNNnxOeQwSNUOZyfrl8fWwWlCll794g9aNqpb5czgFcKxudREp58TKbHcWh9NcLsuIYOXJ0w
zwX7TXLO/ARfg2fUHuBWZF8+9Yg1v/WmhwF8F9IzIDAKLqVDAlZSdKxEziUp+OLOUlps0zMG47nm
F3VbEBIXfVmK50L2gws+GY5n9IeOADqahR2Q5/ca/ciYXN68UA0Tq/+oUGhVDqhD3QEPz1VCeRXA
xlSm6dK+94S5cozAG30yT0fjF+5d3F5wa4IgABLhuhwLCCuR6zniV/IfmDes1FkOilLtC7Ze1QBZ
Ixq5sKNaZ7oFl4sw76wuRTjqu7WxPzd77hCPFf+piUDkZvJYZtxO/+IoR99f48+2XtAg8VyTeWAV
nH2gRv9Pzg9HNypaTYh6FwzMVBUbw0sQGDBM1ya6zA8f/kb6sDj+d48GcuPDhrby1cEspOxp4gZy
C4rEFD+weSaDvqC2itSaVY7G8RWWMmb4ftwiQeI3sxjLCbGcBJTyJ6cRSI/qDhNa4SAfOZ85Ov/w
KZh6/mCsEAxTYqGm9wghcXLSwKpVbZEalQpMg2/G3nsXPGrcT58eH9wLQbMHbh6YYFCl0qMYjLVa
O2A0lUyt4Z/+EKmZOdu/ykLMOVAIpgXeoVHKRGyv1LeysRrju4KHKpgMymqp/4ZGP6NjHSmJnduc
sBY+65cxOWWltN3xXhJEhpqem0b4xhDR2IA4ZGia5ylCqngXR49OUvCSRzKF2PueG3YvZK5wSrzU
OhSbCXWgayG18/JvmGpDLfogDh65NPZOl3nEQ+4xssCmN+AYrtk0ajQ0BwKM/LB3lUZ6lRMdOXRJ
mgZRbn6U53tEBVO2c0t0FZcqZsNzkG/bI2uqTcpwpLtvYIQGCxItzRKl4qBl/8WmNc2maGexDnJ1
4UoiJ7zF3OxWOXCoaXujRtmVi5RRfpUVwVgSNngzpyiIBbdNK1VhzSjKzh3LWEACYOnWuWakJmqA
qppa11PKx/Plw/QjMkhJWVGX3Fn2xDLjVMfrJsYrREBX99junhcMMbzoSngMQFREKT/8/uDykEAO
z0zd/Kc07Z3G9Mv1LWxBxh+DxjO1ws9dSJQhdUETsRwN+aYuFD8rq00X9Sfjc7qg6uYyMIV8LCdo
/t783Os4iGrJ56bP1Ams++SLKkZOtGPoo1jpMs7m3kkg5AbAPjtAM4Xw+tfEKSL2PkDGYelWUqX0
ET+G9cwKQi32TDXyX0nrskrvzRP8uZQGi35ymT/V/OrPiP+LYVDnyvmLd/Cjr3t7Uj7m36WIOL2h
+uDef49tVKwpqK3XYR7VarAIGQcIqXkkyt1iohwYyyww4yBAXCdfexy7AEmTff8Iuc9QhxZ/BEV8
UVlj/l/k5j7yUsmIZXScTN0AnvWcE1BkVm1gMv2rwYEea5Bley4yV2iE/Qzf9MhR0eE+yTxSKr0T
i/oEOYzbbiWFIEjdvrkIbkEYCOYEYbidke2pjUkR33AWHbTrWD8SXyptIaEQ6Gnt4BtzsTE1A7m0
iSaOhpXxY8NjBvbDBRYqkeezm12B+3ng/CKJ2T+U5RTy7NGYtqRledr/X4WKig86I+bH3huArXRr
Lc+2/X9cEyut6klpfdXg7SVmlRdLmfTD703G99HnR/dGFzRrB0aF9ONqYzCzKpH/sECeF7J+9I1F
BsB0yVrPLX4QwjdboOQuXzujQiWlgMTAYzDILBkLUlzOk65S8hxKbopnZ4GkTLXPapYD1Ev626kh
Arb5jN4oqGU+lbqUF72hnpR9lJvPXeBJEvKnFnSwPXl8kvJDQ2LZ+wxgBiCWd5qTs6y45UFLOWrF
SlXaZr2D3s4i5yiQr18LpuGDQvS5KqaZ/typ+7Ex46nHIBX0AOjUHwCoq4RtlsO3gTDSZRIM2hzk
Bj2XEMnGeT44EDMm+PzySw9hsYjyrtU8PbTlgOvPbkt55v/tFpRza2nNIhYNTLr+rZigYXtTebJ6
FAN1t8aTcJQjE7+dqL9gaQKHdMv2cNNQf6a3F6s1IltiF9YPVz9gV1MO8hWq2ZrFnWOaSRTCH1Om
9a7Vy8yJ8F4mpqwsAewN9UOJ+5Ie638Ub/M+avoq40OlEiUXi0Avn6oMmNFQNHAzwJ/wq8X1wmlL
V+pNgX8a5aOF9+R7HHN/JR6COH9ju3sh9ab2/jrcC85V2Y3gQbngkfQgXEfsdDIA//9Te+hDmXHq
7MC6x3zyDFnUaJ4WtxjbW47dRXVRmm2yhz5pgOOCLif5FPvSTxgjuYdaKTzRkFdQom6RdCQqc8SH
i9jL3dy7gjW6aek5ivkx6OBa/sE9UilYpicAlrhCjFm0qHV4NWj9z2Y10qxiJUhCBfYGr5w8NCf3
UtyGHOPsZkYOiZWQH8/lWrLflWtlMg+WRySeXqvNBMCmH6YI1NNkU8/YtWGK+ffFPTx5PvxDCTZx
Hy3isqwWDQgq97P7HpNHKeXkLTy+fvtoJw3qu4REWDbMaFoWMTUl1Hhabquv9BUWrNPyTdhOxMyM
FbI6H9h0lblCRwgcp3RC2WibmdpLn/yhwbcRpVWMY01nZrg6faOTYDMKSBtY9PWvbNQSQ2AVv2Kg
PFNl3VNVLfrczlFotg2oxyduJg9od6kyQtKVrqR0g+jXx0RjRzT7/d76Q6KBmWq/xy34AgLdiw2L
TlessEdotbfreDMYyr8UBHEiHmSsSQyl6rDAacdLM81s9CWnRhmWOQ18xWuWjzPaLL+QBpm11Yld
GCvTzHeuqR7BMXaGJpg6S6zszk7wB1jtkVYy3faq0dvQkA0L/WxUzpqDVa2BIbR/8dFkLkXY6Tb5
mw3ApDIQ73MQ+YdSLlUBx0t0NUJ74db1o/xu/ertp/EKdKYjUNkRd/izgjr8/7df6ADTyRXpZjRv
2eFSDzVjvM62duKw8yllqyucjeLpKSoVxLvDgr0qwi+9zhCWIwXswmhMrBUj8uBZV6XuHcjKyrmu
8hUljeR3X/81tGHBEb2lmpN+wRI49HXktAv30LZj34/qUDmSIjMhYp0DNDYJL+Yy9uRw92fhGKRH
qC0lgpoYdlvwiSEITyK5SHEl/IqwWGXS/MX7dGiPqPbIb63RkPQGJ4KMrpSGXqCfgZKLTTB4cTeU
hcyCTixRSnHzncgZH5vLkcWfI/bMzhx+zG2N+4/3SQten82t+e/8ASn0mfZpYhAp9Hq2UGLaBex2
gS0ZvjeM2/lGg7J90dpVlffOpb/AkquE4xc0A+Cknfrcn9kPnHhT8i2Ag7/5pEnvs0zperMcsN8g
QLM+XG1FbRTHfrfJASYZHFAHlCylhckrlGaCw/FwjxpDDAU6TOT/ZXv85GW4w3KtUNslAQo64Kk2
B3kNYHHiigpHLRhjj7Ct0Bp++uq0d2FPkmgHvM1vPSdxcZo5+pSMLcJ5NC3JRTgUrEnFk9hpFi/h
Sku75e14AUZDNFwtKrf8iWDkIzHUFxKK4m4ywWONSe++8zUNrHXd+Qo0oFDcbnLLuFO8vwXR2TRk
SoooP2NJd86a63lurLjhfAZkiTRENKRe8bSHrXyn07dJqAbCLF+xAq9xq0FfMs7C0zOA4eGMnocz
1d6LoNckSdJrGUn43iPD8Vr6Ev5PdLBAdCwuZr/4QnI8EsRbJpHdgpMkNmVtUT/gk0l+ir2WXPfG
uKZt/covsa8aDR0pSskQdcrK0dK3p4GLMzSPwtnttrA9S7CditTYftcE1l/kwBFQdakrR2IBukma
03nItIbjNiMGYvKnCkcIc6BJhjaMHkdRetfc4HpQDotbysxQiNy5mJkl++vERvyhg1g3Ll2mvvme
meIBzI/2ii079soKGc0b9VyHopkJx+Y4xcr50EtJ7CuCyhSb4coYl0r96NYgg+reLV0/tUPZiHd8
V+yxOX/RaYsVeTN60eKT91u7HoGka4QtxzNvaODea97wQvVHmxZGbs7RI9v9jrO8wG9oidjvvpmX
uKgYbVa7NOoUNnAButgMmoSPMnGkLq3FLmvZZYwajY660+oQu4M1NvO0zIunmIQRbkMNAw2PBbgm
lA86d6aSIpmmg+msks9rohxBp/ctULVEG56STsDfFBIrb+LKLhkBs9OW/Oe1FH72O8i1cR1H4RNm
g/RMsCx0Xw0l8d5g7SB4ly3q64StuC/I9KMsgfB3SgAhq0Wai0I0T2KyX7r90at3Cfq216S9Wz5K
rew+dcr5Sh+Yn4tKlRsc483e2X5tMraHT+0QoAwEZ9yT3TqvuJCcyo+uaHMvF1ziAQ3MgfLnhXkw
rjuoS8qH1ZaLmCsscAjyJj5xcQQq1026qU4FHsBlohlBMiULVLD4Oe6xVwGJOH4kdUp7TgDHAT47
1BAJdnPh2AuSQ5ELpTowruUhUnkTPddcrbkOsBbbQgj5zy8RyKlRcBzpUOh9pGKlU+qCOdv4hO+5
q90tA0Ob4o13m4kcxrogPp+LYqPceUWD1gH8zUbEasbLN16eu61GegFYCkxiEihtUeLeMkg42c16
95rojuSKVu9pj9OfLpCB6ZR6qkOjyjQkEf6ZWrtIsUCD4m+MInRlmgXKkbv6RqVvah4s9mJosu7T
H7xu+2A2ZGlgZVPEJMlPjRGjlCYZFSzkqonGrP2QXNSArTTgKhkvVCz00EizwNzTxfGenCUkD6Rx
zxsBDtRRGRdGfaRBkSDbPgHvKL9E8iSuImu12MiqznYbIUcr3rcGdaKkSww34+eWWupfDBdkgryR
xawuFDHHmG7ilgB+yG/ctuWa1EKrvp1nlL++cpH5I2tHvWjo27YfyzX4jbA0GcjA1NtoUVE3skwn
9T+F/L/9BBcNfg1kCyWE16MJlmQYvLX8BpAb9wDxDGal8x6zZxdHpUsgvhUuL1cQJoML1CQ00JBV
HqRHRoq3s9+hXK4CUXlfRM+UxU951qTzBcdLfkTnshPITe5bepmsxAUiXrdCAKM3ZOc9KKwqcdek
b4in0/2FUoutztpJK9ZEVA02312f1qOkQ2mgn1R61rzu17l3YsYZW3h7o3nzEEJciYhpRVPw7/0B
VB9MP70XwJP8hY7+qB6SZ1vfz8t53mfi/yBRVcUWq2Bc/XZu3RS0kyc2HdHC2rOsfRXp/CIyBi5n
oH9dvVghRqwUd4+/fuuOhEUQPLZqzDXJ9XSl8itrFU0i4FRXTp5IsCBwjhgVSsez6Ks5Dduzebw/
X7gUKm7kGkMss5ZraAoBNB3HMgzpbqNtBY6Fcn3Cm9Juo89gHvD0VhtDzB8a52Wy8P/yP5QpUfpG
sLcXlYqZgDvQcV0EtffkNpYjg+iEbEy8sW3zoPLE4zT/p847FNB2zMGzwSid4R6463KgoOInf0wh
dBUQzPb1sgLfcu2Ar7ggQoOsD3xUYVoccF7JHzL1Ig9BRYX0y8uHBBPeDUEDLyrJ/tzfiseaWL6h
WYNSChEqguvTGrrRlOcftPgKYWSzIKUfJTdcO021yZ8LMeqndpEGleIHdNGUDrOBpnwvmJszAFtf
qjOIVxUe9ysHfDSWKYTLFtrg3EwpsggYFFaCvDiuJJpAGTpKgbWvSB9V5eIv+nDpnu7NX4jy/Wic
2F5xAacu+UrLDxhFaXLXMSrxq3xofrvIDkTEGkxKaBjW7qeRCYZppjafoZjlJgsUzFXfFj13VlkV
kwbwLZUOmM4u5yXNuxyN9TJxoadJvqZMG4s6C6Ep7MWQmuF5coxXapOeJBtpYaU5z7QY4yS1R8Ca
l7PJ4ylJPixY5VOwTF7stMQ7uU6dDH3g+jYxJg2gvX8QtKDlhK8JOts/Zc7R/DJ6qrBVFJKoYMiA
5F0+0Vc8UbG8THgY2VjeABvLsy3GTIuo1jnZN8PK/rADedoDIndr8EMNYfm/E+GgyupwYgq+pu91
1D1Yq4YM0CzGX80mozz4DEiQyE6vSnMRtGt5vfRZt8IczIU0YcVNrGQPBwfEM6lBVDujj1sniTCV
rctLvTzvfEi2WKV1toUeyCQlVu9AA2u33eKpKcaSo8nEwoiWLYTcLpizJT4BxJdf9+h7ht42GuoR
K79xmpgKGnhLeCHtMjOPezZtBjr2yGbjQ8QmU9zBJ2QJBVAeLpn0l1eF+ZlC/fdg+tzYnc+W+/UG
bNUCjddEJdcX5vRdv0JFKAMFnb0VkFSgHv/YollR3K9+i3lWkQtIgVMuWWdehiMPV8hlXHhrdMcD
E4m7Duf6COmSLg2PnSWKLOBrMh6lsBLDydjkeLwsogFGRdAXOACRZWZhqEY1QZEvGk5mVctnvoZh
FxHlfVy2E4smSfs/lYmYj+zk9b2Cz36dI+z4MePbFzDXlvH98iC1BYDdliRRhVF9J9n1qODtrilD
5vUAVQQ0FF7u7HKYtQd0Ryo3tyv/J+uCBPrnf/xtZKvrgwvAN4hV4Ardrvd2Z+kTqKDRYwoAO4LO
L8Sn3Vc47yfFEmsOvWo6QulXL35GA2cKyXgB3+i+nVKoGh4nV6Y6ts3ysol7rgZGftv4t0AqSYya
sGTxoFz6GNDinHs0WPZajLUtY2ji1cYpql1uje//jVdkFvgqsXVDcDSsiUkcTCrVXKtuQ7ANpqAZ
mxJMmkTtdfTAo26Wy/zizmMLSxDamU1ebvqXi4ZB2cNpIwJbsl60jrAL/5Hg2XocUoZyS2QTrC2J
0Zb89uMEW26vJ8aVDUQOzsxDoODqN7GdjWtIcBkD2ajdvjbv9k2XuYLGmzeY6fuxGMnBy61u5EvK
QUNdKmoWcAXMFVL13pz76RZRMXufp6iiXUZQIt+tLW2qD/p2v5KZtCxduJ/PIx0DoxnYOFK96t/b
bhTHUo738KF7YQOx5Plnqcq9CBRl5U8QfYq9uZp54xhYX3CuicmQvz/abBO873e06FZaTEp5nYdX
DhH0RP7zl7+UYzQaxtgtK9TLfR0Fw1oZeI0if/9wd4q22p0qFCG9sjXGVrvnoJMka/yoOP2jY7Uk
Ha7WWtjHy3FGtOZA7Mq67C6K/a5GkPb/2qZZ6Gj8lk6l9+SBCW0zuP4NmRq51x9Hg9bch3cEXbCd
9xA4eQWFjoLXTjG26SLo6EGwLNhfSf5v04DxpCm2NuU5o6AziCreZ7j4Xcq8wQxUdNpJYVPxz9KN
kmbaMKwNvV87I4O7Slitp5D5NKazCXH/T5N/gJuVcdvM4D4o+ac0nbApaCx0TuppyztS4jo3EKOc
zbpQ7DkIYORS1aXKD27xy9MRlCuygE9yr8vuCSDhsbCvswSwKl554LUyNvDhFwHrCXVfDk9Iu8el
p+trNPgZXl7zu7jB+BhznBReC+LjSGThZZwnfopQMjX4t5z5TUL1yz+Wk8+CA16wZT972at467MO
Y/7aVFXev0tKWdzQI5JIRL4NN47OL7FeyIcUf+cTc9u8XUt4/Xh26hpURLeJWhFVXGZR492YCwnY
FgayVaZmbk91sm6ErdcQ4h6SLo0NePomX4O98eQY0yCFOK86UvLvUJWuoWLuOl4JuMThujkerNGx
Bb/cwo1WAu97TS5rEqTG5qwM5F40x7wzZJcTcQolAMcvO+x3lIx6cNHdNdmFlFogWRS632fCcr4L
f9YmYboNR6zVDekEToI6TbwjyenmbOggMkYrVTAPOPZD+Lmx4ZY76OdO4sjlxxSxo8Vjolzl5mEN
4Lmp1bK7QLdXzqMNQ7WW0IZwFDX4GsYL91EJ9/QdfJLi+EKrfSGGraIjIqFajoI2/Lr00XNmJMpi
0QDj/oip2j6nkfDJY7AuJH0mPqRbh3alaWLBdFPt/UjMCVOyFMB1urQlKtIl3QpUTC+TaeEL4Qfz
9sZnQlIBE5ScNG7hLeDefJv2M8mc7KpdzTxKE/oYmpXKYsvBVIt32iaExMicXQSxgbnoYLElGOr8
dajESOF3jwhPLQ1uEgWvdsQoV67aMOSpza7/ZvcmfTGR0nmWvpD9TRs47UWIbkBYQ9CANT/VNesB
0O3G90hzfO+coYiVcb2jS/XKXWM0fcJ+yboMP+xzJvcRLW7JoyGktjkAXqP3MwdwrcvWfTW8H8b7
+dZmTBTvTXSFundLJeadE9oC6oZ1TrGZRDXFli0EDlWKiZr8j2ZWdWi0MoCFaEQ+PEITZa754QET
CphAIK3TFQBYmhGfsastw2givq1EcCm7ADTqZYb6zE89Jp4qNdc4AUy5ImRDxWtssSqajfm+vdV0
/WGvq6cml3W3+aRji8ga1JFPvNCLHOA48/jM9lpD5VqsKaWPRp3/AKEjNEd5zVGe/yarcBvad41c
Tc17p18kIIjsz5U2Wde98jR/mjJNDe/y+VLFPzFPZ/tu9iNJkOj/lYRGF+DUA1Y7hLvqLSuadGf0
mXQdjcanjHeKFDiDufAK7INsDAQWf3/rIXCAXP92NLoZUGNDRI0P7NcUi+5dxFbvXRJbsN+SN94z
7dlBYshJ0pHlY1SVyEMzi+QRXYK5u+hQVDqrAuIMZmwQOi+2yFTKTyjQQ2oWECU54L+/e2fWR+Bk
1DQL4m4QgI9uk/mWAyTM+2CExV48ageSkfwERa/qkugnW7MVyVhN0TzKUQcja2FYjSaYIxneCQS2
G7zgHrbtIpl3HkFANFZMW4IgQc6BMfYTAJtswUuON/QHL/NiPaGx+bbG9SVVYnlzjVa/K6q6vDS0
S7etpRu23jN1a9IExOXx/CE9fUHolTrUDvqcZnRgI/Gb7UmEOEMCOxP6XlQJhROWuLtcavPcgTYV
dME/qO7PZvbBmAZDhi0Gd7hBzIqsDWdGyvVd7jZBGzbA+hYVTXp1sQRcvSo08Nuj7Kl9FhmJ6Kyv
QGOM9L85pvMvWhHSii7XZZmiKusI5J3+Vk3GWopl2s42ORBQmhF+s5r270D1aJfJUC/NSuv1f2Za
G008FMFDYrSan60xZicc5oSin9qQtzYmMCRnoNG+4jWM77Zta6NVmPxJn7TP4JX91onVpi+wTBo2
j0qMZKtFwcSLl0VNpsp5Kn/S6gTFCB1x/9TqkROLNk7tHKW5TElZtOxicbIvOfwabzlepBPQMggT
rtQcBe1MonYwlRqv+vUC7yv3HvXfBSKqOG+clfrT2NBXUq/J/SlfC8/trIa21pLKxSrw1nULMEI4
/61/EzM0OSQngDnVh7kU+XbTFaGGAYVcFfIg+RTfJQZnMyv7Y3iJcK7ATWrcGCzRwJ/NlSlcP8VN
dgllzmjC7XSbGUd13EWNvaxikeMpk7aClVhclVDwf7cSi2DQolgh/x9a8LRTXVGgVsJSQxGDG6AM
GleLLT9P6BY3JBnKOt4/7vuk/24P2gE3zV0wNVvJtbgp7S+uCHKjVKYDiY54oG6MmXjDVyYVakM5
NDLOMLgPdAC0hLx8SnOzZtwVfmtx3eeKqJ4H6ZW9WgVWqMzygpVb/X1bI+BIrxlbDf+O7uGFDu3M
8F6t9WLzRWqm+s1vId/SHMUETAZyni7Y5Tg/s+qcCUcvuYr+PO6PBcTVvSga6drV18KWSCm3OdFs
vEVnvZKmFSxEVyQ0dNqRV2hv8WZn7GypNi7a6pjExVXhfZglBDsi1M518zJHaWisPJ7pzPip8Hz0
I1vKarwxURTBrDCM2i7phi2a+qAxvyed/bmi/ersoql4R/7CTHPOLXUcFQZmMUkJOErJhatz3kjT
pjpKIJWCeXgLmt+vhOVPpCvFwKaGTmIqGn7oCkBAgSTjD0b1Zpe0qLIzgEY/4XAKtO6w5p/L6hXQ
vHf8fkd5Fziaj6azz2tbsQKzqw88zox2x6ifFckJ8TZdtbue4M5hPTvOVdlE2OB2n+ziyRlcHjDs
8beoR2XG2LLcBmHbrgmfmqQLkm57mtvTlfHm42AEl3UnLvUL7rGmmJ7xwPoNYCPz4jtGvGLkCNzB
rAPtY/Yymroh6iAbbpZ6HDiqr+N9YuVhwLmOZ/RaU64E+Re9wKt4keZzvX0Y+D0eV+U/K1PagLhA
t3R8ZnAyG7t8bYavDfLfy/CkfgKBPXD6jINbZBYNkR+PrttviEGAmn//+YH6z2Sy7euJZh/WfE4N
rIqBUUb15Kr2UlW/t7x/HeinmeKGuOzpFj7ji1neyrV89Faw8N4lf6dr266MbGP39SfWIBOpVnM9
ZUh3ZrqZLP0GBUMavL80yBcC1IfOD8erP5GXCPvvtCsqXC/XVYfr1YQjPY2bGMq+rRUTVFYw64Jc
1lJTPFAu4jAj5A+F6knHgK6bVDnUB2XEqUspPAdeJttK916VvxYvSsm3xw1kRrinkgypDUqwIvOE
O2Uc56hoJjWrSy4HojSs8miCtLhBrq7wQacgE5NVq5jUO5B73mQ3KsqLsBv3GQWNOmcjne3SI0wi
aOxm+qjHMBMBbWC45I7CqIbwTdYJShb8UMSomzkBAx+zj/BToEoJSYV9TR+t9t5lhBzQHT3XXqXl
wElb+UcshcxuDoeHV5Sa/bjLmSPihx280IaltkkE1abrvCH+S07Zbrwt7lnsWtfFu+YiAZAl0Rtr
lMMkaAcJJXauYkAOB4Krht6xM+8rMEA6gMBPIPz4ha4IXEyCO38npixy+kvwoOBsS6x60KYJFRkZ
4A0YlX2Pc7xeMyfsB2TkzDMOdowpatBFplo0l0K1N6W/yQ4uVNj+K4BqF/IsZbxZlKwUtZMK4foE
fXYUvRKQeCBNN/ZK5tPjnO/j4eQnO5+flreIvjITG6ZOGGhS340mhqrlMOuHc0XP0zNCCmV78eC6
lM+xrWMWhQb3QBQHW1qkRJb9weXqGpwkiGk+iWpNgyb2oX8mh9/KN59UoKcDwJyJHVLmZb7QuOqQ
zXeU1ZNWmm64vZ2iWOblgEfM/zUCMjbCACepmlqsECcnpjKwljxWWhZ468Mda04I9w/JH86ilKck
WVjQ+oI9MdEDZQiKqjg8gXUxX1DweOsKVnLfmAwSqN/0GWWvJNca2bqFZaFfipSciMUogRMEfczH
OfyUoxFp5GKg1jt4J77ZCjWlsBNDhRZdVTLuV97zXFbx5KG38w7YiNTh5oTMpKiot+pOWrX4aqh+
Y1gXjpVFD93D6Iuh3yOtSfi+UJX78+gdEs5Ft4vpqxUByf8l830wvcMCTjONBHjhY55TopGTrCaZ
1nDY1e/TWnKcyvl93Rb7BrKucMpLir1ADvbO/lvJOYuf1z1op2s8sUpF+yKrcp2PeJqjJqBRFI63
0WiMM/nQr+g6y1zr7sv6ru0nHCcYf/oD6jNtfelCdLIfJmueEZLOEKO1tOO38iOtrlgCNsMxVVyG
Ko0ZbhYo5EE3kJV0cPN6XE+NUl5DZLKnKv5TeaNNHaerZ9FVIzYPFX2wQckXKj42+4q/qS/Uq7ZA
X0DJKgylaMYw/+dKBgyvs4G6JxvcZheY+1BnZX84i/aV93LHujDCfGabfEUUYIyqwxH+7J1YOWHq
WHkXKJPr8Us2kPWk7aKITPmGK7zvmCqTkBvDE8BoYeAA7kvR1IEz95aGHeM2tCMeFRDzGoMdefcE
U8T5mTbck/Jjprh1yLq6iPWVf05mGgpBGdQg6I6n3oXu2ZUEJtVylfedOC7lNqc8u+ru48Pe51ID
QV9oMUV4XWr6REfwFOw+h4Hj3qMixfzj7ESazC/6G3aPlo7skIqSinWdMeqG3g8mHS7s2bPmOZjY
hMD385NEhyCrSIUAAKkNNydEgzY8ToLJjNrh28Z8zCpsx93Vr869LQDJ9c1YKGlYREIU3Oq5co3b
1h/T0+OQNwSikseFLwubV50gjsR4S44W/iVvTrsEmZZnd6pP3l7RCXBtD1ora2ewFJUHUJpgMiJU
HPxVEGw5lVFlnGlwryyipLIJFPbLdzjTq1ewgH9a2Gi1U2rbXMDidepsSc9IpCjWRXt7t/TYh0Sl
bQhID0HSVo2uZPYKu9YNGfcE2L087OS/lYDZ3VDC2tg9czXbgaCXaDcTRWFGH7ayFZOKl24XW47s
0QoGwDPUR9u48VEJhLGvXQ5/1iLotiQdCvyoMm8xlTLAIzjjQAGcjfB/LyK3itpTC0FtT4K2WEew
Ehyk5hazBEaZry7PuSmvF7J4sS/JrGzBdpbb9xRAL57GioKdfEOY8sQ506g4ms8JcjDZ6y702iBW
nZXcjMg5Nl7wooYJZr25lptZJ4rmRm3pEmHCfz/HDRWCFx2gAnEInJ9AFB4iwXAnpX2xf8YsH4Q7
ZQoTUt45KjzmXKOS9BxvSBCvdyaIRo7dmGr5esqxjW1CkYuOetV9zR9ZELF/JPUsCrMW4XEwZMYX
k4FOB3eC9UfPYMUwg7GY+VbMbUX2CxZkoc/kE+Wj7qJZbZtYBTxdQVxJN7xJfXoxgQCPjOskbk84
T7u8HowfyOhv7njNhuDTiOHkmAe38bX3vOx/EZ53nBQg9Ys3rrbzV++NSFyaFOqZCSWXB0T0gCEy
r4iAG++xER9K81r/chNt7KIwfFuVYhqy2CyS9wHWL+/aLR3vjG6GHbklAaZ41MCeweH71UPyl361
RAFRCIaQRYa669Nxgvo91mkqp2DTAF3IuQimY1mCGvuaCMpq9M/Y8n4quKqcNzPFvRfzHupa7PHc
zIYVf6akXgWTdXbN7Cae1mv/T4SOtAUsK2CIQB1IglpWlUdMBg8P3O9seDpmME2/g2tA7ot8k5LQ
YPZM4P9J1gRk2PXtmZxN0LLhO/lzn9CVM2o2qU67yd1OjC1xG8qpqYlP0du+MuzqNOrw4857AF6k
M2QoAtuFCo3AK0qfVfzVeov5dp/1MjwZKSw+Tod6Y3PQCFjYZOSyJhCRpIrQGhcfV6AigHazG749
xdAXxjCZOB5eUrqy8j1mVJpzAz1/ext3kfMD+VS+5NvAzGjI4MXPH495T1WYZX2tQ4rdOCQMVBXM
73P9Ypl27XadFwKEjNNwJlmjYSePaUEbzyaEB3YlXt+diKHvr67d0MDQjSPUJairJeoeEXx/lbbd
8JZ7JrKdVA5+sdTpLP6lghsGex/2/U4sHJZn9lbyjJwXAzPD0lSAXM0wN+tj0nXj5d2er2MSivBX
omHCUAXakoSiN3EtiGI8jqGDfyMZw5QnNu7Bfq8meBnoTnhygdK15/gxfzIVCSnJ+jS4RyyxeTUL
WpNTYX69BXEK6ikotQ+94oeOeT7vO6vrbtMKUqpfxIknRPa9v3ZMVcvHrORSsCXojiNKjwNcY01m
ejkOfdZb6fvQr5bT007Aa20nojqU4CjD0bIQhfTRgEGFGf+rqxqSgnLzaVcp+4g+WoHDZoFOddZK
bepl/qaYiexK6idXNybPCj364B7ON9k/gBaimDuuuuzhO7o+KR60GIsFqr6BX3SS+rZetYxIXhX9
tJywmrHy7WytXuOH3aVuz5N6EHTxgMyIWHNw8mw9udx3A/6auHyEs588hMevYSI3/xB4FqKoOYiu
5d9AYlLJUEQa1Gi7D7428fRe1wtakJVkqZD1CNosEF8tZGCPPjW3xlnLXlHbGV3uKdVxtipvChm7
14G3aikLzqH29AS4gVNlH0HAbm+L+fpuF7BWwEZNvYA9nnJ3v7s0AhdYMa2F8WejR16xB/e3PLlo
uM55W+KCNQMgEeRK0x3MEePixKW4Plw/qFb/LkLFNEJ1O/Ll4Zl2WeBz6kZ2qNjWsALmrj4rFt/7
9c4zQ3OOeJSPEKeMB7bp3LaYLaZRiWuWXu2FiCL/FYUP7ptnx2Omro40gK+7TA7GkLgbOpYaDMPx
E4Yi3TYhuSLe3iwXRY8NTtIT0bIt7UjTTe8MB3Sri60RZBAJEe+DhV7yUpoXSrpt13vdvh9iPBQf
7vPvpg/W6SLMO+oJUqcAmyyLEQp7j8677rk20DgN8gQoyMGpNCvoEAq0qanHs4gfQUpz2fI+yNum
GfUfO5akgMvoMx/fb4B015soTru9/c7fV+RSFn3eXwq0Sv2J5rAOYc7dbjf2ov0fON0FykzeHf5R
bBb5zxq8qQVjm9DiZXJN0Pdka4XXHVvnHJuB05qj9USq0uIwKd+ihTB3edeMrPs19MKCJFGYn4DI
6nrDhU3SrK6EI/YHRdCveSI3szGpH+RF2n0c4THqEP3+lWCkL7MPaX7eGRF/iHxj7CK+52rD8Ham
3Kob2Q7OHm/p4+at/+bkiPx/FQYQbTo7CCIzTjrLbxgF3Zwz0RGB5KQLg21U3U0p6FnGC4BZW0hC
6oSHgN0w/2nMfLvVxJRtLzvJm837mzukHKtkDSbhn49Q69VW9geKXXS3v+VtZ6jLAim7yjlylFFq
sQoco7/k3pyIqt2MYANUfpuiNds1zNtCK4ZsJ7R0jcYyeaprmUjsCeXfmlMNWmbkW30GoGOlnZPB
OmMNmWt/KNgjOXs1HeKo0q/14HWjSsdVAe4RXQK1zSyOJPK4/2XETwB4MYIrt1TQf9qflMmLnNoh
I4LkwXghlLM81uKvdpLXHdtVx7REPEtH2tD+bY4V469QZ/aGKpDH9scf0uckFI44F5KaA2pnyv/b
uYe19P5iADWb8+VsK7LFXmlaeED7HHKWTiA75gbU4yxfb4ixbEh4Yco0KuZMs8XESM2DIZI78o2d
lU+W1vHua9U957DvqIkUFyDeXCub7RuGCudNRMi+VnNaqTeAavmYJk3QRWLfLk/6P6+6JUPp+wb0
VLvE5FSDGrWKabNfId8KUtn2YWULjMQzieJK9FPO4qQLnFscp1t76oo/SHHEkBZG/WmiiDRksCxn
IeVDsJ6Wp6RRR48nDwwtR9wqW4sMjQmfkwRk891T4hoGZIa8x+XPTbXaGySHnc8vU3lB33nmqOA8
RAm32O9QzQ9joO5oR3f0pMbg5epUIo9EBBFEv4DGl/zBcjRMpqDaUhWpz/uqAe+udfJo63d7nJCj
5WDnPknZXyG/z12mgzR01kLi+H+un80p0A33yDUYYmbmVWsFGyg54cR6659ox7xveONITTgofQWf
z39kiKKhkl4kUKHFafI4wemVkjRXdu2Nsdl6+6wd8fZHZ3vx4xMHWC9YZCtiEe/NOPRyr26faKGL
Q1V9DOWd2rqVE3TE7fCbskbycuF+kt6Oz4iV9Eo/RAomwCifR6oBTX3APX/afWIwj6L2ZIAvNo7Y
F7SmvMEStM2Zq+vj9Ic7ZiuBoJEqe6fWcRukTsRoSC6Gp81JrHJ1uF9ZbzWfvsfXWF5t247Pv5C4
YW0QOdtr0QwMHhxgC9JTAy3phVSoMuA+s4fFgstTCfUDREpt1B6kfdkLMWdJyDxQA/ymc4NmGdkD
44phI94K0Lv2H934nmfROeyxdoHufifbo5BRLzPKhTk4xh3/ajLgCbSzCsbgWBZiHW47K2Z+F/2k
YigsPnMfWi6oXkyy6ykt7Wa50e++cAoFwFGL//OWB+cLqh74ggIGRK2h80YMu8M8zpUFprMc/Vjj
Qso47WRjKSR0YoD19dYxJllKyjoRfUejl1FTkeY/tXZ2dUxj7v52T3cC3bb025uWj0ExEmnOi+R0
SbMOngfwg5w6xniVKSZQPH2zPkMjx7yw14Rg+we8i3KyED2iyD0Uy4fCYF+7CUJWuVy3Qos5mX3j
MDpbA3/Ynk+FYSjWLvBU9+JFfQCjAHikyIv3ZJTNEdVzkb8WM4wNBW8xLVMCwTZ2Him+qShZjLMq
OqENBifLYUSeZoBGpNVW83LGfTosEjMO5a1uzebNvjdNCVT/6yCyXmu7ote1SV5t5N2JPkt7LeFZ
K/kFMhmAYzqLxV0NeSkpV2Ir4oCI7VxFYBVpDYqFHNAx6BXrUNyQ1P4/AQZFKuucsbe3PKPyT6TI
WkrHmZfchcaDsc780obBtfqB8qxuNU+xMyV+W1JZI69VwlJ/+WwGtZsKr8WCVKmEU4yfIQyb3FBp
kfFOl58HfglzwD0KvZmOBoNNH7/Ndtksn0YGw0uRZFVByx3jtfZjvE2ACyUCg6MMiwmXo+d7OXmD
5/FPbqsNjKTguac5dWfmlc/3r5RsjYPihw8vfYXs+cq4r4jJLVkzBQd3EXMmzx09eaUoZ/JuTMMB
bdztHh3/ziaqvIc3x9O/XBZ2p8BaOJiGqql/cw8uZRBdscyfWyCMW4S8LTXsVdGo6wRzk5nwWvRi
jQZl3oaiXEC3WNCh+NuSHF90OSLKECSDeesIxADKHo/ZZagAUz1r5gAUCZunjJGZZdVT1q2V9b6w
2cpcauPBALIFPvzYi7zOIau9Gy+YjLK8jfVmkpMvby5J81Q/PYkFSjRDczab7kgiI8sMXsyqwzDz
vhrK0ikum162mmipRKB7YjSsjPP56kTcEcXNMmPRG4R8YIEHAVL0yRj60IQHF3O07P17Lc0LlyiP
cLYU98WlkMWo6QfPR5FkRXwDWdn1ELVrJ6vpL9b42GT5GudmQYbwO5cOaVXvbWCHuFr3LZubS4Bh
pRO+Em/R2mPmTHTuXIvfglUexnl64ZezQEGvlpE56MiSuQiLM12bf7PB2Pn+EYEV5QhZ1GvAHTiW
AqqL5VnnccV+VA2IToBqeYlHOO+kZ8vQn+u4ozCC4qjpihZT8i4cOs7wd/UjfOm9gRaOuSF63Zp8
a99ln1p+EgnMNTm3hIbjlzju38aPJBUrlYeV0+htqAvwOhfs7e/cW26JA9QcovWUIuVnrfopusV1
wBUZNdl6drnhteRVilghqrwIDaC1fxTDxtSDC8lwxycxzzwI8Q/pxkeTxpZltoBAlJqJaoUUgN8I
bqwtxRJn+ku0+hyDN91QmSCWBa1pccFcmI8GKg3wPfj34pBP2/9G73tvP3NDHEcEHaQLS3wkumNy
ZauXnVZlgtMRIe8T2N9gnydYUkypnQTM6pP5TqMHwOl/ozj/+u/88bWviuwltNIkav8mo6VlbbUy
H+0HNHvsBwajvAl8Bb3pmrOs/ZAdaX7lyiCIjUEPOoTarNkyMAdjZp7pYfF2N+C1JRcU2wTMYqiE
Ek3fzgbceBxbyPdqYq9iyC80AqpZ3Haj9bSJbfy0kzxF6Gv1MHH7sIFNiJD2zyeUlnZlYcj/paoD
DcpMHQD6CcHM3g4Qtqhq0EukTdudGg8HmuDmtNpsLRIE6kuvDiGq0PSPDG1Xj5KnYWXY9+YIW/8C
bJI3wLG8KuYbUKJttG9B2wq+iWIZi1kqUJKEwpDsfmH5msLUG69kfl38J+Kj17k7toob2NWIjjxQ
dIHQ12RmAT+kZ+ZFhxudy9XaSFCV8oK8YnZvSaFa5fVz9a0oKNIgX/5Jq1USr9+Am7Mklu1c1wSV
kRoi0ds7qJN7oCB/PhuiMCIOce1qooKe7VKOTbu/r17iGzoPwlHfy9gEf2Ip1quV3n9Q+4LOq4fX
inHXasCTRkT8yLmhLzT/UBaUW7EcTd3aKv1Vw/C5wWdHKKhc/5Uyx9CL0u10fDKQIuaujephlfrZ
Uj9vxGr4SjqcAX2CuLenG5jfzLe6tlpQLrZqYZXwbe4Nw3+m78uo4DiY/SDooi6yoB3ZZFVXQk+G
UfR+1az7WX+YJ5CjI6QYI6Je/dmrL9C0AVZdRFf+NWMuxGE0VgTaOSab4Tmith3JPX3m+MKmuy9B
v4Nk+Q6EpLML2+cGz+ft5rse/Rp4Aepa/BtoXKP0VbeVqeQtvWzjaDtEhrLqE5x8QP3XZ39gMVSs
WnUk9SIYCGiLOW/J36Pf5jk3E8BiQ01vcgOBSbXQeuM2Qusd3FVk4I7ib9rL00HYVMU7qGCIP26d
Tf2U/eh3pUxNVt3CzCZdTpELEu2MgdA34QIUAOp1my4Sz3A6a5A6O9xGzztxy9yzj4MHh+ieACow
MlJ5fLGCNDN1AZWfVHn9d/Lc0KxXZwwKI1KCCbdACwB4YYZfgx2mCm/RbKyI9W5UTi+8KXyuoQWY
QoiRqs6u192tSq49JvvjIuSeG+V+UsHsqumPkComxlcLOSvXCPKhPTDs8VpIxi9kbR+phq6wL4VS
INd9ZTU1hBDJE9TcA5sTmrkJlIyd/ArfTEn576fax9rmhGyMkS83XxZo/C979st8ptw9oK16zDEP
XklNS9YNtTx7lRlkzBlGlZyJCp4uesduNCSGGpASmSPSPbpXBO3uQRYyc66bDCKCs2qljH9d1upE
6k0mhQVTue+tYNo9zRDrPiAWsCZnJ63/mfKGy/Ztl0fc8tyBbBqlWiCvTcG3ndV3sM+unDM6G/Q4
xJxHyTzqLMUitZ8I0TZCTPi8kJvJDbYlXyqDQ6hN678HGpQn2TMF6s5fCmk5OASUdvu/ebxD9LAC
AZwY56miwCPbi4baPAkaS10norf2PUFu36+08J5ALASiP+voCPyt9Gzhngm/rOQl4WMIg3ZSyVe1
5GhLp1efTLp3rweAIo6qOGc58+K8tS7P8z9foVrXvWIc8QEiiaXSGG/+jZhTinleghrTdPETjX+F
btS0R2NkSnpi5Xyjieu7eE2LbirHPp7GCxXGnFrk2Ip/kMDRxg/YKdm64bDI8Li6eD43udWsTqlK
79LMG9zYD+GX1WtIZ0Spx+ciOJ/It3gC4FKpYP6Rs7rNNN4vbG6mf6NZX+V8X3Trh6AIORfmHLdz
xal5YrI410PYVK2UBQXAv37kH+QRyxlvibeEv/nx8n76ZhWS+GIBz7gpOo51Brk8LghxgROX0Ogz
9DV7odq0u8T21havyaAlMwRALovUOR9r2o5ClmOPP1SF+U1cwjkT95A1MHHRTE8okSguEA0lVbSt
gMdJzNf8ZM0VqnAbK84xyXI6+jyRHDDhqySbRiRWjG4ZQL8EM7RvVM/oQA2yunPUMf48qQ6rKWUz
8NNnVvNlqvz/ajZOhaFmFk1djDj5P/Eqq+D1spDjdmt46Fc4CzYhjptpDCxDS/EurGQYw0wEpoDb
59ynMQ5uinGVRKVHCGNV7S6VHOXXJwigd3qdFf+O8cJO0EWWgcER/TQ0NM0cbHTfsPhcTimNEwtp
vr0Nv1gL6W9z8atVCQcBfSZbD+zkeC1jm/BU0YI6McrGlu63JbFY16W4jfjo1jS3eWFhJzJUTIkf
70th1ZAUFfAqSvQK18kvp3Ko/+E5873pnHFvzx4Rf8U7Pkc4OPJZfxZfklh4O48bu6pW9nXY3wNT
qm9taMmcQbuANPGohVmIoyKakZNzE4aWymIZUJ9lDGqqgGPFXMsto7zjF1q6FS5vz4xD8MLp3jf5
qTPiKVnz+kUzQ/qf6nHX68jfD1HuC+JQcYxKI7haHlnN+kw1ELrbb0CCbqg1SoL/BW6CUm2vxrnj
HboJYJC5hOD5KVTvekwpEM9GHQOxjr6qWKaaDbSlhpjf0s6c7Mn/0/1q7DWa24dbEukV3YWoLLdn
qKUdQH0j9M4VPexIBershjOPixQm4LuqFy3v5RXSHQozokRW7Mg4GRIvfX0B8qJLi5CkOOZ/O9En
JshBDO4A+zVkmRoENqBP39dcWVEmHmN53Xm/Z8yomMQ8oyu/YRw7e3yWnJz+DuB/JqjXZ7LlhtdH
aW5WuIzI7sGg8n8c6utLK/+Zv5ylouZ5877KD6/36ea7pbv+iigoiXczqbcjgtohjlLitoL1ZXoS
HvgkeJVh0LJHMMx7MBFmD3FsY36i4aiFemxLw/Y67UP7PcDYu2K+aUgyH66cEhoGGSGfIkEXeU89
e9rLRo/a9lA/4H22NNJhj2ML+cTdFdsukoHBySo8mpSmqvtpgQDwCzpCfNMIvL2UnncUNcCbaZj3
rrCeCzqprnlMgXsW37/RLaGjGeWOkEO1bNbWphtqmn/oS3IA9CIIFs6zXk5FCqtw5+ChCPEVcqzJ
zn5adoMXuJvCkGA8g6Bbmliy4fD9BR1o2iIuAsXc9wBn/wsn20IBEbCZnpJfMQRAIF55eeMQ8qbl
RYREoUadfgGJ989JNMvHk0jqcbdgQIQA9Vk2g7y7k6wK0efYVzff+loFIUQuEGONLmZevCufMSpg
WwTG3j8w7jboezf5zGE0H6C94xHpD9W64S9sOg0MSbTbWGpkCpqCyMHfEGfcWFY6q79rtcrRUdkO
RDVI/DbnIKzIs0F8H04RoiRKgPTh/1ydcdhMgtYKUHMH+jYyEIcDvkbrLEoVcouAhSP7kj3yJ610
t4jvKILdjc83VuCaSvR1oexhhbhC7RvuBgGMTOHoqJ9LUBek2IODHJ2a8EmdW6Nz3zqTcxmqjQjD
6n3Qti8h+H777qfhzmINJw5fYFFZcvzPz9dfB7Y+BySzVRnR+L8dmLy0r/Wg62H7+5Gyzyhgi/lq
oCf56xqFkNd7K8QLspHulNyCJrNleJIUSkBTo51W0s/MHXeiNo9MdUBM1OXp21CxBrSbHA/BOJe0
HBXX/itZsRS9/jwnyPbgadNJJ2toIwtPpvCrsLOphRjx4oMXlhFUb5f5bxiamMDoZgHZwU8dMnTn
R8XWpqbX6SR7/UAQWW7DxbBzeUWDmqBhRXZOqH9mj3Jf//9ux/PJ2eSgz/VFtY5FvabNXCE9cEoL
/JS7URY5F+UpxlC9tV1UXYOUGFREV0HhDf3I2DJCrhOoBxgfKobE6SJnnRksH28sRZ5RnJRxFH9R
jqbXEMmz42kPwcOTiIQJc8ZoxVI+9220rrzyV/y28bhJWR3I3EhuofMpfnROazMmGbSSaT+9KhbP
h/nm9zncwQAa1PKi3DrwNsbtqUSCTEK+almz6+Kj1gcX9F+3rmNQUr4/hsiQPCm7KejcEnlmppGz
2ygxHQlKL1eXNFbYCa09JWU2UyT74b3r1DFL0em/JX3hh+0IDUX3YYRsaoafhM+BUvfNJqRfGocB
Fma7fGgFohHRmS5Yfv/AKzbYea9s1ifk3p3gZWEsy8Qr3bSple3nWv27xc9mP8HnT+a5P8/KfDnX
caR1XvGrtQyLSdplmF3Qis6nyAQJTZ8cXY7Tx0SQZhjHMfRtU0a0qPZJvEMZckWRD6CCXWzEAHb6
TL23Z4QoOYk+j3yfxvU1BOLseoUGpz4qomMHEnPnCMK3VIRzt91kSm5NYoCg+PrMenO4O5UoYAnb
Hugzy4gaI6yWuH2L40Zo2+v1rjRHnLNgfFTd4ljg3qbMktrPn4505iJQmGW0iQKLhCug8VcUvXB6
mMuSb5k7tw7BWNmD8WAU76AdT2UCi2ouf6+gbq4xr/cfD0PkjW6Zq6KIY50w6KRSyQNU5Rv7yPq7
V09WlzwuhNhk42wi39LN5O2cEq1Mf4Yc+TKkKK+YVUItaKcsRXlaewJweViCeFq2w0zur3LmT5SS
5m51jIqGibTWP9cd8hQMGrW/55/RoEzvR5HF1oG/K8ei/IAZFPDj09lFIC1R+fSCQ5aFYgq3aFbw
cHfR9uNkzKHSEgewhTtkk7GC/Ze2J0qsrBsJCCHg4vrCebMUMiBBJLlLQ9mN9+Qr0DVHJyen5zj/
nPg3dX0FaOVIWvhbWQEMGjU8t6alSFSnhx4ErG+Inbymq0tygyCQ0jb5Ty/V02pHp+QfO5mkEmU5
ulI8XBiuErgYCM7+1Ci65MwcFpZLRzI2i2j11XudBOMKaZrac/318vMTRKDbgQqz9pIzHAiTDLs0
ovIFVCkuS0lwewkMqNoDHmNuh+E86KW7CKnxQL/jAyPKkU5DpRdmp0HTypu/7qeCu3ctEgQprvML
2HWypTCq657z95EXCLDRgwYb3K1JRZjo7Di7Cko7SdkZRLDNKQpxr3CaTiYI3brMsHT4fHRIs4Lb
DxbkczI19Qsjnnfg0SYIR6bTESllNurE6JlEOusQzWMbncbjyQ4n+n8ovD/mEZT0veKujz9NLPed
gwRAjYA48Otj20JXZJMvKi3itG7g8h3wXwnbPfhRnUDaPnjtChjkbjYvG+RhrPxe1MJy+7wAqubA
U9MiwLH5GAdi/3SLonCI5wB+8DM6DSIHECMqAIcjI0YqzrHnpUGNrHWfWPqlhUOOUunKKRAxw/+f
26RDJBe6Aa/3L75oOFpatCE4eDhY84wswH0asZz2L3j1s2RpR6B+1Xi5csGrdfItwjD61iEUT4dt
f37Q4FnJM2mCPuubfvML19ASVXNeUyFMMK04hGwwDJJk7DdVmIQ4nMjKEZS3mu0f1OE+emJGTF7R
iwrj+RyHqdj44Y6izU6AZVs5zIip02Wz2VIkGO0qlijCZfxtcZZu7HG0b0WBnvUlKNV+V7+5WoDy
I/l821c230vdy7XZF1DNGkJoXKRQGD4mQ7mlgqlRJoJV0OJvdJzpyzTcmiJdIDxdqhwGFnT5g/C9
StAm7peoy6v5yWeWqBLiTAbetuXVXalnhQ7QnY8DwERnohxM461TYNQCnAFtcC6N+r1yYawGLaWo
f+8S0EcVKZ28ZgKKDr6b2+8hiG9S+qYR0FqcO/sc9Blx6e8+vP1ys0+h6W0fOK98vzCxVPQ7DS5K
x10US6lccdQ0Ww1vHymwxL4TO1A32by9Y1DB62zF4ayEPQKJYCeTnCKM6CXu3NcNEsOYMNCSGHVN
W4msJgbf5m+PkIcdVkZl/IfFoFydQSQ6eanNCsght6HWWBGOaeBRQefyHmTWdSsp1ttFsaufd8dJ
XPD/RbFIZHcmeSOUd+Kl/MWwl22FeLs+yhL0b09WjlWtIGoYXnvc+EsHCsrmKwRiQ6vlEpvlK6Qd
BZOslDzIP1r4yIsZP+eDHGZSlNu9cqWsdLmMbea9QtXRtkOa04K3wL5QOArYZ6EXi4de72VKmEF0
cYkOu6vvd6WcqLy1X6sf9G3cEFO2yOtnVSlk87DM1uiunmcrj2pIeGnnpivwsGoOzuQtFfEi+XYn
RD1WbBY/JdKCW0IhnzseX9wAVwLJT9CnQksuqiIP89NSTg1UcGqFmmZKGpY2AJOFwIegdsflJUEu
omPRjA58PjJ3X5ufw6MffEJk4nX3l7tWKqsqwA5cD7gjKzMzwekbWANFY+9l/fNHbu28E6rgEl7R
/wtblPi8AfwHvLyimYCAfhcvqhZXonOmep+R/FCwl/i0V0zEgjsmY7eYl9fgzL7IyFLz73ovTWJv
4f76fgACo5HIQTXl/3afQrP1R2d/F/vW8Rp66rdrpZ4gWDDZz7wk1sg36M0iQk3KJhADTALCSEoL
q7xDjlk16CezOEiwvEHRF4eco4lc/R4NVbVTJ4B+HrQlpJtb0q/vNpkd8PucP1TRCg1fWjJoAHKt
KAw3z0cVnU/LdZSKvfHQJu+ryuhOLotHfoDj/N8wUpLoM1KVKp+UqGmlOCT+VBuOWoxqYzwi8IzH
wJ1ruTyEk0d3KsXZzsDEQDKGUON7J+M+X9+8jgfch07362tBhTxkhnXj4eHcUm7Fut8Y0jGyFZxc
GRCPV6O353qspqhgO2RIpm3+jxc1ZcXb7NSt9UlrSyxmXG0Nk++kvXJ+S2rocPqzKqw0BRXmBNNo
d3H/17cWv7xVjszEMhRL60e12POHxxcYTyV2kPaXG6quzsHoZ7unNVOjuCYm7v1IMpitaMq+9AOp
ZUsDqYotXqiarPmOKYfG0Cb5nPeFZeNjwXQOTVCS3noXSj6xR6mjbLzBCQ1IZ7PpKGwCjh3C0MyW
Zp50WOuiUJfxV9A4Z/kH3ilhcSSCagEWDLmj7/Mo/3VhW9JCv8HqcK9F+Fg7AZxc5skd+qQjXnuS
sJAQxqPLYsm9+QgkwL/6HPCDMcknQHvPqyPvT0hF4S8+NyqPvOIQMd96Mg+CWu72RuLWLUg9buR6
lyC5ULdCtvvo9YoNnHmgtudASX6SoOrtOySB9GN6UkPMtHNWZPUMWOq5XqE8ZQQzrAvuU6npdtyN
QV0mSNaNe8u8r7ZiMx6gQGrjB7BvL7DWjbfZU039KXvCwtJBfoE+xOHg7zCPji8te4qky63wgCjN
XDmAulQ+Jh9UjauLl2/+2L3MNKz+tmS0T+/6kwKHqMfph+3Bs+HF0czXYcaFylq7IhmiCTtJlBL/
i5yMJ8z21tHRSJZMthDOG244H28WFO7Gq373khNCOivt3LOhuhn7COfmZXJJuMJi+ersHK1Lj7T2
kiX0flIUEbGGPaKGGgE5xm5wkqDCxujEkomVOQ5gjrXDETQ6bQdeS9vFYKZ4iED8feC0De8guur3
yxPYXOwbQ+VmGOE6P16d+4kGGe7AxAxPd2BkBuCS/z5TIQqMeq83DZonYRwH/ih/WerK6tHGzxlo
l/+w8bnzoVF26gzQYMdlWKWi19peWat3T2ZBp4dOzlU46BjhccR5BdeBrqoNArIz9v7uujoI4GFW
nHq1fIl8GlK2D2vfZtZT9O2FNKh+2zAEPi3Hv9mg7YYQz8MEGsY/3nxNsgbv8CylpQrjl53r+/Ig
3IzwjDKRn7noa1N65tqONvtBLAsgp9K+jWbteA1wsAOsp2AJxLN6Xfi3UYsNIuYsoQndA2Ln4zN8
xR8SEtwhI4TYPu7q1aXkeIQ3lMv6ONx4C9Sul1pWpvS9jR9FXBTzLKVbxWz6hFgnt1+Dpd2jZ6Xs
y8Pho5EYM6z4VKqlKeCghwvfx7YzTHq3Imkvz3NjfE6dLamWB3wzRtODYZ4vAM081n6prWWBYoGB
ftHRTCrpxZuRysfl/kL3YeQibAUTvnRijYN9bHOSEPR2Hd/05ZxOiAgmjSUj/AA3ARR9gN10A6PC
9ybNIXz1XKLd5wZJM8kGaAEyv5TMbQ1yzXCugB/AuDSzO1hvz3o8UgeULsN87NHca2edJszwn7wx
9/DMTw7Vz9mFrxs0lo/E0PoND64lg9Sg9aea0+lFmn3DcMCAoJNcGw19DGFE7MNJN+wXOBkLBvqH
dNtjl1Vs/+ezE6HXQ/4PN2cn22aZ/hguC6gV2pF/qCCb8T5SdRuGlBfkYt0z8TN2Gwtwsanoh+Mm
wTxLuglFkCRvNPlVmBMfiiLRieaYxlUgTyUmuT6Te2B5XEJhqxUborHUjow5tvRuSYVlqM+LZrVX
hEYpK5HmbXMmIX4XAG4WH9IOc8U/SA4/Qy0X3+eQGqvpNn+Ir0ar3EoVIdG4wCXB9VJLYY4sdhEe
9cWd43A1wS30OS5s+/k5XIH7HQHw9U9bXgeuFUCvuu7EtKpWMSnwXBzZX6KxKnLH+7lOK9lqt9jt
i7Y1mMBpno0/N5sCd3zh9YbqyjpUxTkmBF9Sop2IRr79fvbfYkBt8r6hj+M2PW7+XPM3lfjOyacV
vdgvEXsM9JbrovtEwqmA3Goxg/Lxh4RKksGtb91XCYHcjU1KzcrXiRjafypQ/xZ99TeYH/BDeX6T
kevnY3BQY96ctg89AILyAZmpkC8h3Uyeaw5V3H2YYuqv+adO21edsQGok8d0HdN+ZMKHGAnU1HJZ
b2xBcs+wvmHohgEm6YGzkip2ZeEWep6EXEGBRzfr6OyfGbNOruwL9mAQnk1unTpyLgsX/uEQD4cE
X68m/0B9kdm90IYY1AsGxR7iNJCx9dNmJFg0ANTfPmxtpGdYHrUe8bOOOYGi+OHx1z4H4DBUQHJC
xxnqVMT9RU9C6eKtq+EGtJsS9Bb34xP2vFVMkJXB+zN2cSqkMglDjkwx6XL1F8q95hOzQiD+4BwY
xntcakpaQ/vSpEaC94JCdA1PTIwXes+LLZXZ2O1mcIlrC0PY8y68rD9YCW9xmwXnHNhHgAATYsha
lz+tioQvMEJThCMGY9TVWjnNrMrTVOvW9faCFaby1F41gl8xwZriXFRja67aUQs82RpPVdpohHTW
MePQxZj1rlSnUqmD77SXuLRmdOWejXGALOrk2Dq3KiWCdhiAPer+huzFvwraBoXGUvDOMh1AVDjJ
eftyI//mrkgBLFm5EyAgBrwrF4U+r7GcThxcAh/1FG52GJyw1KD2zNJW9hkuARVsw++JLIky9IYX
f+xI+CWFs0VhBHukwBaPKp3DIDGuUzAtqiN5siftp5O6gfX4wJ9NNhV335ImBsmEYyRF9tlw1wd/
BCe4+LFFSSsU+jiWeR4ifTbSXKdBgN8IM2WXJL2Lxjf/bfru8o4UEkSNxNtUVrkiT9EeVGmUzbuw
BuEn2NACJXXhrjal2gMoMzwRvuCBXdejwiBE5nJNtiD0OY2jecCHiTPHY0p8cTI5KASjy8kM3+b6
XWliI61uXlI2Jl19wut0uzudUD9l9iEDv/tP665nSMrMENln+eqAF4VDi+0LwXdhDHOJg8WHmG7c
Og6rvOsEkOn/ijqbkwSP90nW/8/bW9IOYwHfVtFUyWPcEk722g/ObmavaWA3Jt61irhhufw1Ioy4
XmBH9rvwl/m5VbI8xuv4DSJBypnJMaS0Gn9zfREtrMWRVWj4ZHawL53zgxHx2LumULY4r6w+jigp
2JrUcwN7CISiPKGZo5zFl/kE1RZ0w8FLAYeCM9SesCoIypbOmnsZNZ1JlbVE37/AshD3HS9zevvV
EVxXBp/khuAJ6zJSn949eCvNvXSsq1ZUT/OfSOiktb5UromcHfqjUitP97Ri4fMZepJkPGejyiPi
thLkw3Cyt1KoiZA+hHsoS9MXJFf57LglAGm1zlqY1F5uG9bWdDwuEtlYpS+C532jAoh4SK5vmwPD
sBYCzYL2mXRpVE3yq16zMY1BspffFhcpouLITKySL85dPA6pNDdDLQ0zXJl7ZKpV4iZJCOv2OpTg
WfKL6iaU+2hgvC8ppK/cuKrSs2tYRbk5UgYq1bMRUu8dtVSmgm+mGPj1FIVdmlRX1Vfc3KRdNgQS
1G14J1+6lYiWCYPaEvrth7qzjwDKIDnlp/AYIQgU0FOyNLQcy7RhYQRTPQ57mtcah4svI5irQjr0
d99agd05t2mSEk33/MfhzHNw2LTJ5kaFQbxK99YHagynrFU8REKvpzm31ap3rAQZLX0t6IAHn0lF
UiHXkdxnrky3KvRsOt71WVbIpNkiRsXuyKV79tZ9ajkkNqODIfhkTGRyrFn0+4M41f6XNLN6SrFp
16cDNOfHgPyZpT7oYw9uXEMaPe6u4iEmLVOmr5TlJ69z32i8CN4Pq+oEM27/PeCs2QrqtJEP2aOf
e73DUQDl6FHN2qX9VvHcooong099liy9XQLUijfYFM8vvKhT7qYAERsJiWc4ndgtSKPg/U92laGJ
Yjp9DKbWyVLhFz5vi8RflnW7Q+okriHfwclovbFCMw2D4Y3R5q1ew5vTG+UoRr+VZwSNQyXfEEt7
OIVkdf8BOMx0hDksjGxPhSBs6XEdpL+1LUdTn74q35/KaxYpgj8fdKODEIr4QyJHlJgn0x2Y1aoq
fibu3iwCnGbgfNWqEXK99T2hS4+3XoakBB7vsj8Zvmz8YrEZS3EPdCn7Hjzzct3go/uddaWq0tAd
rds9/421kMAQzEYtfi1RyHcp8S/eHLjjVL1YtmBvx5HnLfa1WmRU0920tyNHZ3gcw/wltB8y3RLA
PyTibhAKsmPHVarsQV8EIV/Ngte/cvzvSqIT5PYZkt3O/AUcPJKxRE8RLvJzeRi6qQqUukQ0XtId
JHEjS01gTqpmMF0RUdG983x1ueuoxuwGJxeA+sDalNc3FCXIEG5NxGZ8NJdRGL05p/J2UqgMXFks
B/c5Zj7geqZhkouHsCQtZJzI1uYKLKnMUPlZ2Jcx/NqVCzhTKSgV36NZPBlCJQSnY/2jJbuKwYuj
LYtMLgKsbnVpzGt+088ekVp+/Ss6Yg5upM+FPHLlrmeRlhX/2GkjBqxNQP403baApMToOo7WAdcF
o5FQb3OxQPq4sbg3YjiIN3TCsUB110bfuRbeXO+oitU78yMMvmFJsB3yufMMWTbiW/PJXvLTO3KQ
b5MknRXA02VDRYQfKsHRMfVI2HIuG7Qbua1cNp92cjuxIHqcygQqf3O3ZLj7gUNSiJd1W8QmOLfy
uRIib2ExXbrfnBW23vt6gFo8Fhwd4oKVWoFiTxeRUjH7rTjAgppGGBR22ApZFV4c32Zvt+qhQ25Y
2t2nZnpF8eLUvp/V+tIdasrC8hErRqc6KaWqLXkzEK1X3rCur/BqevcSPu8ZDR7gSpoyJkNamWJS
aaIZc1XG4rfy5RwbO2ojXKBkPiuBovHqjnBG9A93e5KeXMuGra1cUAHQJyRfpi2sHeAN27PRlWCZ
9kIz9yt7II2Mg+jeQ+23Sa7/K5m4ukIQg6IMmmWCsyAs+ztl2cbcb9D9xRbkWvWm5uAjavmYeBFm
MCiwMFSRodEibIpmwCLVwhimorJIWsYxRbXUNhaAtygjJtXtovx17IAsKeGGviZMwvKC1USwNLEE
09nrPfnmZlcWy7nmp3HsSi4wCVu7Ok0MlfYGHj2VJ1jPybkqckEick8vNhIPZXHPYUgJ50EdTThW
ScU3TftJMkfdo1NZOo8hepawUzNSbgo2iLbGLFk/m1AP3wIn/d0bqLDTWMOy/AbKN3qpnLTS/Ken
qIasikmN2ZYKXIFYPwSx1fP6OdXDslhMe5h2j9ut2XFbuTQhb1CBVN1uMGSCtJaKvSgyvTX4LKuE
cBuFd/hnJPY1zkJkYR8cK7ECzUx1N8Q5ADtpws3vw+RIF8s2mSqg1A7kIfwqTjS+0GF/VwCzr3m3
XFs6jiOvA+YbnIdPYvvotTilnG4RHmOv7Lu7KZFoaeBmyG0xsXnQCoczuNBdDBcKUlvG3zgM1u5+
aqplTodXpvn3le36B3PQW4Iwm5/xzBlMJvocVzrLuAdUwBZVMyMVRTZPbVZYk6kgLO/PNh4fiB5b
H9IcIAYCxJT4NopQKuv2MTMBRQN7T/xbaG42iA7FaZ8Jazw+OLZuHN9ROwaQeK1vc043T3ZntRfW
nP0DrQkbPN2+JkhT4FQ4hTHlOD5Jggn1Ej9bW4TYPcYGDXPE4xRzOeqFBB4Ka/0nk0fU45/WsNAV
AFgDDt0d0CKApq/prasLB/hs8eZLfk+uE/jx5yzr3yFyq4uxG4ebvjX+K+H7nHFtCUsRKyPP5iI8
DGpSRXWrFgNToOpdrrpfKsCgt6oKINZQtpXndauwZx6lr4ez9WSdO7K1qzCY+gEj1iCVYOSw2bxX
biBqfHjQQdpTQWupUvxpVjEDY+uFZoRhSUYw4G3XUZ7RROY4vFp+flWUbeAxCI5gS0s8hdG3rO6i
731z5Gjk/FQmAZ6XeNI7dBYLhvT8xzBcTuowwGW0iZ2wxdHiPk1bGJPkmQfwksifT2xWZmp6Xr5f
LOVMCK5SRcGvX+8Y+BylfYR/q9V1ZOp91FyH0aD/ScyxWUSXXJ3bGNCv4u5gdv2TrWl2133vsvOU
x2U06SIT6ayQocySxsSPlMPHI4NJrFyxK1IugxrYftzn9YPoyqy1mIEbXJZsmwwPcZmoLNnkZdmF
72MjVj02u4z1F0Gnl0OYGtnO69lK8/leFt6aAUVuefVGunQ/oHNsSu8j/W7lwDjHFDUDi2EE0YRq
ez2OAjVHVg31Fr3rA9vRseVfoQ3Ob1i+jnauR+Jn4uEDjVRGsj5sFLWiVNQ/OPWVtcwn8Ojgsl5G
0PvMM7nPIROpAWPgGXcLJvsL4ieTGSHCbmLtO9lGTcto0KAUxsj5v9gywFSSe5kYbNzG1M7cSGan
p1o7eLKqyUHjV6EgCtTglUvGerrdB2NAa/HGtuS1E6/Z2Y20HJ83BaMxJQl30r/c/9WGyiy2GK5N
vBHeZvSB5ozjwZhZolMCQMHBLDgMmeB5ryDCuZt1G53UfAyx4NgzJDTSk1dN/NMswZG0UpehaGpl
PWsMonTKmBHQbjtwlhlGbJZT+JoUi6dscuWtKDLmgWmYu6ZBySlsGS9SNzH2uiiwTQGqorjZPEvR
1SzLsXtlxTduUUpjMNolaxlTG2aC59T5O0pF6z9sSNa3zPM1cZNjfVBbYipPMcNYkVKuLNnhpzAH
WrTiLwgsnPETkiG55FMZGWA2IMQhK+aAezC5tWAYOu9FgZzVQoHIl93/5ZGdLxWDwnh9wPNIjY1v
zSXBQ/JEwIVNxmlShwWj73EjkE3YsHfgWWoIjPOUiblSmEydlC+raysdr0t49JJXWP5vWUX1K346
CklfcgXIvT1iKaYsWBfbit/5lSCsMQoMm3nQ+0cKWBkNInMeuNMWH2E1CZfvS77Sopvr14LI0zh3
A8DhpGsrPLIdZ5CdApvVnd0hXN+/kXqte+WPjkCqkNh7WxAJxIU4XOHT3dlSvDbW8lhYxrlF0284
6JiJH1QSZQHl0K4B+hSODf1IwnzXkxDE0BvFoo+/e4f5Q2gs5nCSd1SCte4tZqvHb/CQ4F8eyUXB
6MPOjs3DAQgUwA4MIXrtxqh71rEK5TGjbiMOtNtyKmmfRJvYnv7D5JV196ztn1FlqSJEIT0rrElW
euPa44m5PLkvXV/XVujldvFDeLG45rV82f6ScXp+vKPPN2/2D1PHBmBtSQlHYjVNZfqh1PzUC6uF
zZK4Msj+jDjB86fSaCi1QSB1O9QZj0/KWRdGx2treDWQRv0lfBqzApCz97e/8bWK4HwSjKDOEwF6
Na1WSjl5Yf6rFWQSLT74BdqUgdCL83LX58QekKH706RPzBuYITbZsBWk/caXXjcP1NMcfb7wiYjb
crDRaK98YlRXvqrY40QFfMRy3uo21QHSEpopRVvQwSYXeJy9fXsfbw2FXOhr1Wa1YuZT7+43bR1H
+ICK+N0ZI8lmjrWONm1vfmaNjCi8dkpP+YdPNraCoJ1cxS47SShmA/6R5s0B38f9L4JmEB0jThJ5
tRX6zMCvZsOD1sN55NtkpJN94JurCNWBsf7Q37bOTGrhQ+ExjdA9W4XHNykWtRv2VZz2wb1IGA3E
ThutGb4JqotKWmeo91g+KxPfC5+PWnoSe9ugLQotxp/tvLNQolpTZQw0R2be04H7hXsyeMSMjfNh
6TIpbOkbbSdmY9NNTbYN64F3iuLORC8m5intBVIpkdDC3GbYCROIHh0sKXzWXtgkXrm2kPnpYc3g
LEuObLoYNCMLsmhLBg7LhJfJX1g7+DvxtsGod0HflFcvlYfK3voHWQ3nqrzziBYAKpEKPc1dIFsR
1oGCiroAM6cEP9Jjq9rA3xRJQ9ACtiO3qtAPR97v1Wlmjwo5PlII3bpM9k01kTKiXi9v9CDD1Yjh
0cOCK6HJQnxQtcyUJSwg2a3E9X9rytDKIp8tEDHxcZzIb2mpvsJxdB7pE6aSqyRqT4/Abt0gky73
kIqRN/hYJaVTrzCpD+SAstRKYnFkJS+0nWriytk+GXjHBOC8AVHhCfNBkVsppHrqNMjgglnSGzJh
PFHjnBrqsitgUg5s5godVSbm3bChKa6zs2JX9vSZNipxbwZ861o7tKaG/XIuIa5QImkfYZkBkWoY
smPWA2eDvdzttzOHGqir+UO7Idz0oK8yZAal8oOpOt6CQGfF+m6ulUVx1A/aV+jTzoFE+CXUPEFk
V0x4JolgJs/lC0kDmKd62uh6mtlC56rMAUEtQequy3TYepBAXiyJBcA/PsCA3V7ri50fmg5uFk7Y
Clj2n0uwL7mE5JT9aL1Jhlg3AJgtn4xSG603lJ2uXQLgYssOp1IXftHfsJIbpvqWxfg9sFuftl20
KaawOg6JZ9Q1AAJAjcck+WThVNYn98vT643Mtmtp9jiBcW/Vmx9KlO7DwyfbT2yT7aSLeLg1S01R
C8O5XZ7QvDPFBpZz1jnvmT+7klke2s7Kc0Zbu69rWPB5DMloeG/sqW3EW8U5xf7+RibJOmVMcGt5
kPvH51v3JeX6YwOkwdEiLnZiDL5jTtfN/d0doEhWk32bthJXs89qWqiUPogqgkNvGvToNoruoAuv
4hegnfoieBkKOK6vve55efjnJWMqiSoSmietwcPPRWOKRmJYjy+PWKLK2NYlutcYoFWQ8K7ZNrB+
qNjYnR0MctUwfv9WNL3ex6wsi23Pu3XLB8K/d5gQDZVcEynSypYWq8XV/u+cNuth7kv4R4RGZJC/
S4S9xmfKWbH16lvAuEM9br4R9ue4jdkpofppti2sFRr9wy65mV8Gm8nL/ZOY5xz4MFfcQN/c5vmk
lAp36lBA9tjYWRBU1wwdKREQtIdDHUgGv7ksE9OGzuP7sveAdQD2WpF6oMDS1KIT0HSoCU3jTnhz
FJjZM4f8EdPXwxLeCDOMVOXbU+9UwBh1bGZWWrsTu/s/ZifZyBviDNOWCFTIjs3nrBn2jLZVPIgz
vWr0D9T5wYkL74bc9X+7OtO2YffAZoSAj1gjacUt0DO4TBfDbonLPG9ElZWeqjuIPcawjloAsGOp
NvxlPAihC2O4VloRoj1zEfHZkPyGlX4oQ+h8OX94TFlxgkESwkgGW0xqz3qd+1snKn90Akfs2Dn9
AZIDzrBreeJbWXy1kQSeO0tKXqbjT0laFzAnFIWxfoyd5dDwQ2Hbh3gvr6X87B5FcMMM1tlloBP8
tHSuSEtRD5KXoW2syL9oH6c3hXO6dj+rcdUd/hg8J+MBLtS+5aKpgrYj+0HM2kHFJ4LjNqnWlwXF
+QJMzRrR+BgpSzxVrXBXfcbVrkH7QFYV8W+FoBEVTn1T3GT0AN7dfuqPOY+suqPnmOWeL7ENsu0p
bAv4YjIQa05R82zNNOmJqTU0KOOgi4V4pfkH96zeVUFzyLcUDDS6IfB+LB1mj6yGcBxayz+EU20L
V46QTACz5Br+C2a1s4I4dJyX62ZcXSdy/zHfGIOfH4/yjjH6SJtkCtXiBrnIfTPLjZ4t/Muq1fyP
FwWNf+Py+rhxhxeQ5aSy8fWJNBeEw7YSYTSC7Wffo+Q++hiiuNGoPdyTDyUIGw2SUg6TtIwJSqFN
R3RfkD/nw2EyGdjCfNPnjezG8OObr16NDxNbWDSBgM9WWkF1dJZVZEJanjwJwFcNhb8ub1S7+KZ0
sWpi1rxFqS2L4S8hN6a9vcyGmcUDYPoGrudFnx/yNYfmyz/Bk3vcprwKHrLn+NeO/Z9Bbz4aozl7
uSoUVi98moqoAICTuVzJA4QrCiFeRdDRvwoiduYDxbQwZOxjiSMKVumcWrg/57/nz60a4tEcnNm+
eG1hy94kPZpqZroNF2Ga00OnxPLKQf8gld1rg9+NDEN/a2jdWX0ZK7z9ZJM4P5QcNSWShYC4UPnD
NDnUw0d4z1gFzW8fKjxOrO24UOvOVrUYJNpERefIUoSygTtH9D1UFtE+RMMc9qY4HI7jdCt31sPW
+vTOovqF3NL/TFdkkKTaTunWPQ9c4motfBLSIrYCXtaKSndB2+HkRuYpED5fZw6Df4ds7BLGNLOm
Mwe0hcEn2X6BqGOu697xZStfxltILw6FBR8TpwdD7oEFHOxy+BTQzcmEIzYtAc5D9QiLhhRWysON
ZgU0QWWM1FyMbgtYG9T0nYUEY0t/CV23tVSUl8bFhgYLg6ivEcM9eTd/koO0TDQr7gAJS21sGS91
k9vaaUh1AZkP3bmgIJHM5bHwVk7Uab98kNs1CCFZ0Ax9W6hrNv56tTlIUqEKijx4ixZFdt01Ap34
mU8hCxvt5r6Z7hDGWdyv6TrPmOF/veCCRiePtEFOkARdtkLtpSRzv4CkAs3Jx4t2knje+jEPwdvF
CoEvYXYmdXXFEoTSVjUoHTPwrJp+P3ZsAWdrAeaDKTQpyF85LInQnq32ekbe45BjTV5+D1EXgtWL
uSZ10dfFtVtXYWsOQiE0OfxmQmXbdjflF6Huybotw/yiN5fpQXCxMLLR2BjGO5Y3Rb0DorZ/X7Je
nXXs6u7qCwi0lO2MOuc5jDE1tHeRgyyUPEjv1BZF8jhivRkb9j3uRegK575NslRjOTzBcdVBFuX1
OOV5hnxpbnc9Gw/vRagwp9pGkspLn4/ZrXFgYINNgAbXPX0VLONGWcPR6PKgA3Ho4vdBzuay6dVA
ty6vsIt05hzvd7hnTenjcPUYFzok8BlXmS6rhiREnJB0GpDA1+oYFlcVd1DDDst33qvhTJgEhb/n
+vNeKY1EekB6IIbHOfVKxXRKyxu5yT4lwDFdPNHfHvzDDXFWaHxvYU8KSw7F1YeAvveDRQw+67wU
gNKznHj8f91R54Ew8xLOq+DxH98NB1ArfabzCLPRyHH0JEoBRKIu+nfVUUGU+NU6xp3rJH2y7z5b
1m+GUlDTKfXo1Rl2d32Y2hYEJ9x2lEvljsWzrvm/yRRijvHDtU/dkbbE1IEpo3htPUqV5tsRTP7K
rvas8K0fNIhS006nv+M3I/KjsS2BCnSYioiLFK+uWtxDOI9nI0A6w3RohRVqvGn8LD/OT/USLDfR
6yw9bK8lmMJXYJFzjwO+RaWgMiGXGMTc2NWrq9DJ6m2fBKegD3mxaT/6/k/Grr7HRNaaTL4pC+CS
ZMzvao5EFvvMN7A9DtpvCgOcUtQPhsVC2+ld9AIUFCJ+ldydrUMGfAiAfxb0dZIEYztynlxdHCvC
Cf7QsRKxT1LbzM40dhTx7Z1OK0AYE4prHkds/i1qYHS6EDoCD9HeVjyWFkjK79Es62d3El7xctZH
i4+D7I7VtXgfB4nyo+37jtobPPi5osyvf3S1B/2Mp5t4W7M/ukFQwolZGY9HuN07d23LvQ8rL+pF
+KIi4BJm0VXb1fKusnIZGlhzJvmiCEeY401XV+8+WV469YBo66ylNTEfrGRG+86jumzpeuuGqdz5
pHVF3bZWwGNoXuljeY3pbuF4dL0IL0OzLyy/9gsb3QFRe3zgTp0oo/WpxyMvLlmcl9qqsIp2MuAB
Um9ps6f3snx1nbJfHViSi0sgCfMZQybqHWgAKQ8F8T/aH/BDy71mvfKI6M1ebofrlk2pjzpD9XLB
fOAz2aB28fJ5AUos5gMYc3Tb9BNz9YoR3ds9DYE60Y+axkWz0zjVFRUSpYIMekDN5mW4pT0DRV7E
kmGZkrjPB3XhyhMmqqlsY8jHICTFeQy+XjGS16lbVBqPXJ9lNXrAf9At3cnX4oW8DhiApcNXSzZE
MttvCbR3uhYzQ6vQmiJYg4uzsK4FQJo6WYC+Kv1phpfycEeHXOpxWzGC4eQPWNRX8AX6hz9SUCyk
ipcLPT9TBEHPtanmzzzKWOBJ8pXUZgZ8dkIlUq/L1EGz57iqWZgDANP18P+ohq8KNWLZGKi0LezL
ySPGlEzPjntGn6qfKKDc/5PF8j3RyiXtB+0el5xKdih3sprrN3PhR8bhOMzvMaSbw9zJMXe6V2hL
FcxXhyAr9CvyFkXqbry+fXTUgYE8N6qfko+dh8QhLN2N0dA0om3ShZAbMYiKe7+9qyXEAz7E2JxZ
DgYQqUVBMRZvBqGJ8gsdAFgonnIPGBy9cYJTluIDDBpneCYu7WUs0fSgwVBdDiCw8EdH5HMEJAZO
Nz7SVF6V42AMb+UdCEMt63wsixxSmYtv3wAfmzQvWTVgBc1kXapSuYQ+nVBhWUnYyBvZoHhECFK9
BeC2m2ZEhXKuLgj42tBPSC85QZvCRKnzdx+hAkxxqYqtLcHiExDkoJGIWmOM/DYX/GJCUpMH3Og8
p3PlDcT+bD+zWMWRBid5LLQtjv2MUMxt76qAAngBaaOEkOx/uAByLE1kZW3eGK0b29sMTecvIA7U
IfzCOF3oaw/J43VW/INFEVh4jkhpWFLCqJNtbAWNc1SytAOU30H1OOMTMgrGmtZWis0rhmDXG0LD
mig96iZsGSEcH0xfx0qC3LL/unwkJt9nudlRXvf/r6A72kGMAiU8Huxx4QbtKjDckfGKzI06EmnS
6dShuGjvhGyf0y4fqtBJNEWHg1eedF3Dzhr+FJTWZygbep05WyyYhykfGNtnoD/ysBpH+xMKUJ9G
6wQ6QpdiTvLRLH1NhSuhfMyUVTjTcI1mNmu7i6YEshDD890ihVl385zGe7EyRxMooghEHcQ4YZKV
0AW19ZeYF3hqGSJPWgjwTYMhgM+N07lZ2wfMi7GtVpVX4+c/SbManAQvRkTF8La4xLpGbs1zL/qn
sP7oHPrw/PugQ3zsL2QVLfn3+9wcRtPNsPnTARQflnf0xdkP+Jqi/EGHfc8lnq/P1oKNylVQPqkB
dqyYHYLgST+/eS/7YN+0I/afEoYijeCklPmUHnwTv8xzE/lssBXaC18SunXyFws3m1wRZEHqO6KI
OCS1ZKc7YDmMKfjY1wuymjp63930zAmcDp+T9g4lbVZsmlb3L9VZdcsUx3Y9zq02Ygv7XOWDui82
+p45n5GMgjDnTN+h73Ih2/xqByT/2tmCxK2S7bTzrKYwX7n+2xVZvWsjXCoxCZtJfyIC3uL9cm4h
zVl5J9v0KOPcuB3EJ5yHUrjHAzNQBnXD3NuRqYEProtjRQcL3c4MJvb8OxVGM8mu/VkfKOSZQvM3
2BQUEfxGQlILnKosfHOG0XfuzemIfkKtsEFwiyJ4ZJGAX5iN1pZ3kYdI0K0TgG+hRD/Nx98zkePD
141gFPYGQPdmh8omz2dFnS6DOXslOzIDIht6aPqPWvCI303ZHXA7EEEmGs81eGB3y2i9iaSfl7Qg
wC6aR2m4HB7USl3h1GxSZ2WnCenVrqfvuT/VGYlnWR4mBuAlObfgmuYY710B5BvhrP6hpLuBKTEP
y5+YUQENqgt/h6IN0QLP5wXGvZRN/T1HIdQahnLuGqzZmcbG7tymle4GQx/ShAfQLd52rE+2yPO2
xPvd7LRcrcAHYUjP3AUCxrZfN6gEd8RarRKNdkTBlrbGS2dxJaA3m+51hRKBv1OrOho+dVnpAjDZ
RdvsUvzKovtmFVNfnIRS5PjlcAaSFzIhXiEnRP2Ivjch8WwereMga7F1QD0MacIEC9DocPNWroj9
Jqp34RzzQswMBqYiVefQ3TteZXqyqcw67jRlMk6YDlPI0UoXlJQVtUsuOwLm1S4R5Uhazwux22U+
cbPXYzmoqlo4qfRsOrON1b9HodiB4I0RID8WDSZ+1Qd1ZZm0qj5JjfYW3NaOAKeA7QKWI+zGBXpd
B7B728VMXFhmo/DTc5fnaKfZVW/cKi1jpMDK1MpsrBgEsSkp9sC9BnY0KGxHU7EmP1U9HdzDXmkk
W63VD6JDsv9sGoIgA12rDUV26w8f7VshrXTv4LcP8tl5BMeX64oDtR7wDaAjarDC+nWwsoAN6guO
jQ5RKAtAC0bii638+WGH5KRmyBvMFbNvubnZ22yctsoSHhBxXIS8s5zsd1BDvuxLWnpgfcrYADk+
v8/OtxxQwb3ynzOtmyzoa8bXqIam4zID/8FPTKDfoisXQfiO3okWFqClxzloH3ZoCM+LnX72sxnu
UZm6XAb0YZrbOlaQWnG8DQiInbXT1PGFna5vvX61MDEYGYg6fZ5CQ4ZtyhYPQ91HvQjbODnjeHUN
D8Xz0wju3YaoSMsk1U/X6U6mjulPLE4ncQhMrm3k+9LPjTFNoPNuOVkyGQ8elodqGFg8y3Q3oxqi
kk8Om83CUiOn2RHAtCgGPG8QaFRmQSgQ+vTs+ClQ/yZNx+uvNAaTSdRwoWtxbydkAFuFFLK61trm
HVfT3Ifckkfpoi+bXctkMxy6YNI7aofM4AZ3lABbpxcr4b1Xp0FXWdhBIW1JbOh49WvhauBQ/OZc
zbDACVrDjdHPKK+/HmCSSp6lc1MANgWbkj9DoNegsHHcT3uSIbN/pcZ5kWTp/Bp2Nm0dkSO+dLWs
BruYwowvaIfTQ6QmK89OvKH5QBKSQeU9lp2KYgbZrCfBHr12Pf4dbtUVkbvQe2w3+ReUCNc9eA9S
C8EiHHPQhwGV7+fHn1GDmgqWTUNOvMzlXdHWwhsM+nbbXBvlWm4/a05RWhdNt0x8hnr4//MD12KL
Cg3scFnJnOWZjEDzTOJLIl6Yu90TsU73CdWA0+AS6KuFfKMaMJIXqbN1+oBs7fEXGFiCFoKl/sqG
SkS6LCO7letZ9gcyZOwutZlPTMBDnncOO+LSI12c6u1CjYiJppvYN2VDpU/4w4TllTqkCYizkdb9
dkjR0EKYy1q+xrFh2jkRElIcdfBAuZCDtTxzYXaiUITatqUCfts6ueSmN0EAJ7F6Uj7oJPCzRq//
JHkBCuW4NasBwK4MWpsgACf1zTYOG7/t5mdm51xRpTwXqLIqI3ktUUYo593P7c6OYJ0vrVnuBjmW
4NUYQNBoD9iPpgk0gxC+t31CglhK6HfPRaxfIfwqOxGXUYCnP2Npdi32A/4tgcm6OFz6PyyddFRx
n6ciFpxdnWBl4sTr9GobBf9Mu8RRBZ1ChWzRlKjriWF3tO4uHNCyfOJXB2fmil0dJNgQjbAO5gGJ
CTiuHIfmGpSR2ZEViOw/NTU1Vee5m/jKyl7+LVYvlxWDjyWsPnxgbfebngT8ls5t0WyJ4fUGRekX
6N8Kozf8spiKb+gmCypAyg6L9XYz7LL73BEskHyXe1DNC6sy1fYvGtYbC4lGybuMlhyVf5usxBRZ
/3s/2v8OCLYKqJ14wRtZ5KQvJjJrKZhus1YggJDH7VNBBmQufAG0sWXuaQXxKnYp7Gw52JqGjme7
HfL0Wgs/SlbSuJtmmTFEP2ZAru6hnVc5K9t/3PWUxHsNsP0h0u72/dKby0iO4KHNAzE7AHQeKOea
WrqTBurNNkI1RNz0l8+7mJlWwpbuhzdWB78CR7Wkcw2WS4f7pFxQ05pH/mO/VN9evseOZ4g0I6BC
4guWVB7bWHzzyOBUR1QKh8WLT0Uqnd3MePlyv77i190BukoVtuC87LgwqZyoO6mTkulGWGeuWeBg
S5HMjE3Uvehtvk2LQkLgI2Tvk6epczp/90V6fRdmze2ifoa96xlDpIDXKoE5ZYYCe9GRSwJIHBw7
acPWmEF7lrbQkJ50ZE3Y2bj5sjcCP448wQU81XAqkLnlR7kMvm+Uu5M9iNOfegRqYeE81vscR/0A
47Lqr0uVixxOhdl2Ej0TP0Np7EGOvMM0c3KYPAT8LW69EtaA8kYfmo5ZpVjMqiuhmmi+aDxhh0ua
R+fZ0SID1BWOl2+XF3RXLwXC5YKdjAmKQWKr6tDCtUK4xNrpnWJ7QpiwlPdN7IXakfeTtuzG2+KQ
cavdCNx+QsfGazQkTxOTomTMClv67uzpx1a+JhCOSyT3q6vP/osed0IZ8f2+3QxaRYOUlf4XhuaT
emONaXWI6BzbCETn9QPzsvo2jdBdBSid4YztdKCnPeT04QDR2C0E7TE/GKasMxIqWcvayyB+rcIv
rviGFEYZcT4fqLHR4IIB2GGGlh6GeFXLY1/FtZhIh03umiNeccFVz5ymzrtwY2BNm18ZXWzVlGhl
jIM7jVYwjmbpxsCPJD7FkH9/D1+CAi39Fnlt39t8Vo8vCLk60OHx71t2iEyAiv5iJvZBlkIhJjYk
Ht0QUgxDQJ2xohdXGdtlnIyP+/meDjX2ihztGVCMmNkwoHu2/X9JqviNz4Jbn4GoIAQK2XK4Rqof
Oy8lNOh1ChkYoYjbwMTqhLUneXMtUY7AUHzDLtsWq14l3IsrT1A/bT3jnpXlElE+r1CGJDSekv86
bWoocyWrzd1zUxzNWqx0aUX4HnTmHrEtadoGy6zcaBuECimblvftZ1Hu+B7AFcjr1aEbcd1iee9c
5QcRYonYv1lDtzNYtwEZHYwXeRTIiF4VTpBJ8h0Y4gLH15tklQwreFKtTjGbyu25ndllpOjCJHhr
4zZtFbc+orIWITbY6NIgR2ZwyPJTwZoQX/CKTfwT4KgsojR13i1Pjta+uLUaQbscdlpjtoTody+T
62QLKwwwyNspgtUILkODJ9U3KrBoyrKy4R/kNZ2jpxq+62lU3VLaoIlzU66pGY5D76K9/1lF9vY/
JjH8AfQ76B9VkPkJkzYQd38qMdZwm2PMsmEQmCbrnEg0R7XqhKJkGJ0WGCCbgeyu1derbh1mvBli
2399NR4lU0W9z8AQuUpMk2eVL4t8ISgva+nkYMDtGxZ69GZpWOMoWG7wzDGIb46pvaFn9+SM68x7
vGt/OrECbP5cmGSqxGsFV4ZL3RzXUsxqxrhQbJiC0QcyiKquYQenT2cq/0eBHs6wDFf3nJT/pkaB
/SMHSzeiWjLWM+5UkWNWDkOxW2t/0cY7TnD1YfdeQA+DiSFiaHhexfv/uyWbfIcPvbQRd0hwNlrU
v2M4hPxIjxuT2UMxQxETZlsxVMiOjUtXhRSPqn2naWBfMOAtXCGBRzj8U0+GhdthNOPgT9ClhCKO
rPDuiGkE0WXqqqz/YiCy83c5/tJ11HOsS+9v4Hb1m0qgI8rIh07HpnT9kLfOPkbSm1T61x3MjDD6
wv/0HmnDSrQb6pq59n/YbtuTx39vEBzD7u2a9jJQAFzoJN7U+/E9xeuf46FXCxwDAWJ08jtT3UB8
8pCDFIS9vBW4tJm+Bvh7fqHr6vr+TEQ9hdrGAo0XHK43rMkdRHLXPiYF5ewDk9e9RtYgXdw4u3V7
AKqRC9MZxhvpqeb/qnRXAXYXViTNzKZnLQLnddlHQC50kTSbSOScTVSYj5CNc6b8THAPMB479GdS
9X2Chn0O8pL7b+j+1LbDY5N1eMSOSvm0fIJOkvCazUJ+xMHY3qdeNIckixH8zv96TWEPPWjQCn58
5QTcz5+9xrDz5YeFHt6iIjx84SC1LhzaCmvQkrniJOR5litSKRa5LO6IAkFQaH8jJ1lNCk4woA+A
RXIz5BLw7MccWCI8/TtXO5Fpqt+hi03nArpkqPCH4Z/gbPv/RkBDRzni1eAqsPeo/gxw2DyTMg+C
eeQ5mR7mPcAWKhVdzdFI30ltkN0FBOfWVrxTD91kpmA94JWiZREMEq26VeRkj+ReeJN5zHaAWyZM
PAcwrilleF55fYQ3/ylrR/l2rgie0EfFFrdgfoyLFdul2SXWy5Ic5cj/3sd/YvruOBv+O/ANu1jV
wbqU0K6gxuaSJfFIlRrVHwIp/FSMCP184K4D74NtoDVWse3zHt2UVIPIyE+kv84fpEguiH3f1RBI
Gc0TGCw97scf3HUTxtBWcj1RRZVUjPamATm9gej6ow4KVsX5NX+NW3jl6+lHicoab80gILT7k+6K
lbFWhz84zjL+4b1HQrk+Qrz4OztTWEZ5OiT5gNtQ7/uGt7qS7xOx7LjpiaOZgYdZocBVFLCKtL5t
rnR7cqw0lLiqkt9U0QLFYTDLHsQK4WCnzv2yVK/ijynhYCWmcu4YzWzQL+Bv5ASfHWSptlk2wqTD
rpCVKVUgdWRZctcZt/ixtHhxMB0w8SV22S8zYJmejaNkBZEZ2bueP+D5Hpnn8DHI6Zy+M8xN4F7v
P0oNndKN76bBsmpMWB8rIAjphTPop3E7cllC9qWjN6zHBs4fzu5P6XlhFXXL/nmNIeUSHV0BdXxp
8HeSACfoMM+EX+yjM+7ujq3zxEbAGxfYr5a0jt8JkDZCVm/qa5huURPHOUsVMRV3f8/WdGrmQr+s
qFDJPw2r9o/c7aG1alhZGeWpLypD16zv80IqLtvWLq1255sH4rcrKk1+3OPw/Jxul2FoxOvD3t1S
1Re6ey5pcB+pd7k9pYtXeUwAAEbHi2yevv3jKx8F43egYCuUzhxGb2FE/QqMvZM0gPUftb2W71b1
3COKO851d/6vWFmrNmVHLmKwwkt8tp/Rhhg3kXGAP1uRuFhCZF0CsdctsAePm5AUqpw2jZKTFk0U
QrxbFLyeVIQMKdKsYHfmzpKrXluQ0Ce41EfwRgy5dX4QUwFzmiqv4WZtuS02laUct6Gk1x7vRx37
9pms/beN11uVn6Q4jqPZFDl+Gv6UqYggfBucnrlQ8fqzZIirO6sbluBZiE0muOmujL8qK7cRZ4EL
i+aCVdMFf1h7Oh0spjQewGt76YjM7avoIyRIURCqI61qaVXZQ1yhPyMyqWVF2JLau4zAblepeK2G
9pVABw7/dbr3cVj4oM56BxNiG5eK0VerbvmSf3icFEE95IeF9HTR4nVRpTb4FGJMNfMNohQCs2OW
uixkwWl+DcUtN4T0DukRsJT2hEDjfaK+xfKiDc17kBhm7pWEt2QtFuh7zJ/jntTljbPlaz3h2AQN
3U04smFC4l1Y5xV7bUajJk9CsqVY5hrlJ0g3wt/czYa4XX8zRZSmZ+nnOBqjMsRaPAEQJMcVvxCA
J4XVQwTW5bsITUWpY/80Grs+VnfOih0J9MNcBmIr2sCX8Q5KQrccdL+sfWrLZkckEoBp2n3ZARGW
z4Pazy+UK4kzUJggAH7XLAEKy/36llXGuLlIu/0OCXNo0qRA66huWRggsYbcblnbalFJxbsavvpI
8nUhTBFnWu8w+LfmiMIfZYHWv6NRJ7HwN1PE3KwRqRTHSnYqKBdQdFSakx/0VLYpr0owQiwQmUAH
aHR2kviQrKGFaNjpOyouL73vhoug7ah7pb2GEpm6i9n2ZQBlpAe7W0S8FvHM7aUxkaCH+h14k3V2
R8QRg4J1ZoyPXIHelWCbUhsqiwmw7oVSXbqHuT/79Ze8Fm4d1xEhKQc6lAnYm0xmTMr5qG3aFnvc
QkFba3VUqzgT+qViVpUOh6ztVdAWLJsX21VXLICoMQBKGHgr7OsSIPYyB04H2nS94wuOO197GTSO
pDul5YENzEE7eDZVI6yHC3ks/XOf/+RTBkb+h7s7qqyfO6rI9AOsSH9xLlLVXeEct2tEHYT6+XYD
sz3A4+XIwSB01HfgRVhb8blmplo5hKF7lfUxbUIDXUmOg1smW5PNloPTIqDTJniNd/r5Rga3c0fV
dKChi3bGZIlcwHXWowTbkh3FifGUnt7266pG1GL6+kYmdXseubEwBhu57Gl3m7L9t02Woj66iXsC
g+IoGujpz5ftQqx6yVB3f0MuOU/NTIZKIbjlJWsIQnHim1NVE+MF2N4VoyYxOUXNLrwaRd5i5IUz
3cNzScm5IaPTj3iUFF7EJbYl1/owc/DZThGerWaZ5L/yCc6wV+uJdXsO1H4gggwXX5iEplMqvbZW
U6LkinlyvUBBv1U9dJV53G//FbPe+e2pOche3DiK9IkxYs0MhRteS2V5J3yCaLbJpeyWm9kXIQPl
RGsj5HItr8C5LiiI9UjBRqhRCyqa9TjVjnxwJHzietHEJkJpcmWCwN9vsKb9sc17XOaw49ZY/4aN
KEexZpbqULxw4FX3pING2uZ2uiRS5LkwQf4GcPuvpT1of+gcaZYVmmDMVue80dAqI02ZYbAG+AGO
ied0wfVw1YrNsfsCZLuYeT2QJ5F9MpzozyTJPuvw8DoWFcJUx6mngE0RFy9JnDqCQ1qIhnFrhTaE
ckbMDp1Nh1+OmZo3V4mWs7ruVR2QDO2+MRtYa3h7Ue2SAVYOCgSaGrg+WN4RHZe2irsKT4a4nCDC
c+r61fupdG/MbnoHGYYPYb2iwfDgve9zW6DLcb1UfkLWHRCKzScy7nT0E4EWNmjqWMO/klEpRdPM
V5f+TlqwE3JIDuoKhBTKTc6faIQyzuuE2GbCACYdEaYepWCx+ZA4nKFgQLrBIBoBQxy2sb+VJXOx
zkbTugKuuI1fyEhu9yIxiT3T9zIhWnR+HgG2boD4iqXbNGpwLdTk3k7XAIEhkwLVe22HrpeY0/pr
khxpewx8mhs31YRpXy5JQO6PcpJJgsCbH8vOIARzuwD6cT/c8FwF5gWwMsNXQQfuynTFDqpukR1/
FQTn6iP/vaZNTii2kf/4FKqm3hoQdz6MJHEwrzqs/nm2aCcYr/YVswR3hK5P6+wSLrFt6XCx2et1
uVxkLkjGh3+17kptx0Elu5wMVSlOQCd3UkgunvyXvIYg2OUC9rS4ccQelMKm/El21dv/9tfMB6IF
YnfnV3zbPsK/ZC9Fth8x+JII/9ct8aL+5CbTdrdkA9Fg56z7g90xsYStYQmlMrDO+c/KA6gHOz4S
kPf8ckf9I/e6zdGd04n1Z/aqfSCcBqUIk/RdcERC1z9maZm2g0uq3VpgkK9n2Numj18YhfWU/l78
xPNlYYeXaniIw7jt7a0PZWF74seYbhYYmFEBMpGohrD+3pC/XoAKHDs/xrm9jRHYJMhMCn8/IXNm
TJH6kdn/Sef5+SNgymhl3YOiZxKohOsr1PhX1HmoAK4FODG2t26oHIeQeRgpjesw73HQjXcykkoT
D6pBpbNFFbpsXiHBkRAIS/miLpG7C1xRWz0Vjh4pcyBAKlY55C4cKmHhFyoeqbM/lIVpBrtxBHey
mO+wmEyrY3jG3tEKIugygQGUoZodq0x2a2gVyT5QGiXLvyTjIMxpK3DrUlDrbxtpKmqE3hbmUxAm
tSsS98bQu05suV1XkofO2BKzvzqCbgjcx/cbD50yTLS2u897k8tcUnMeMxoF1mPV3HoYberU4jxJ
ECYN9CJx5e/veA7H1cDV5q0BTpXM/1lijuNxZl0OSEkTzpx3//KDwThmHdO0suD1rRtZqS0O7Tmj
pWfMCWf90rinetXaPrD7FGurzaDQ90ngo4XI2JsEl/Beuj9ZqcxlfQewC5ywsuRCKxoMOkGFmZNG
fJ9De0QFgu3m2u9TUIX932Fq9/V54sms0/pAhHp1VStHEvSBcCz2WZrKvCepzFl+ztvtiYhIYqXY
ByT2rakgTnSo2/Zm1/1VLaHaBWZUKUX8Avo2a/pERWj0OuWAV7pkIWCJlELGSMRT9VN+AdF92TY2
5fGqwdH4AeBTWrpqYX67X3pUD/MfFjTNqwkf/14uBpmAaEDTdXZKzu4P07inMJExggAHsMlzfGQG
QHHWObpxy/MD9w4WGGzitZVIPM+wJMRujKDce7zk+t3Ua1aqo8Lgi4B7lCeOPUWUf+7wvVTmyc9v
G6YMZkmlp2EUDZWuLbgH6iCJN51oifaON+mVBnVP+zZDsShspUgecS1Pt9D6rJ9a/Yh0rrp/gevg
2MnWrg+vPEaDQrBlGmqqQiTFu9X8wGdI1RsO0yA7CCIXSwL6K5MEqvYEB0T43G4+gIKWviuSJ5d6
Zq9q+Qi3gDoGplkYO9epg0to/xdKgU99dRpq9h0m77/nVBIaeod59YfkA9zdnJENfjJQVFVFUe/p
WgleH4v9HW18sJIYFb9Jof3DjmCUKlivalcZhqxRCTqkGrLOw+9g2pnKdcQUY/LS2uYogRC2AiBy
oJ4HEFQXkfV1dexccq/5cDLp6UCuZrCmShysNAgNLmvhCSaCjvqAD/MRaLc9axyr+pjajRTbQ/fJ
dHYPX4OIO7XRmf3/6fy4p5GUx3ZNk8A3AukwNOhxxji62F4uTr/ApOLYlS03MTaGIiestZeQ006V
9Jcw+P7wwaMiPqKHeqIzbIGJ6PuzbnxLmIb/pR8d99StRT3tuWDXw26xuvmGji73uj03PatljoWc
Xkna8aKJQOKSlJbaAy99Sc0hVhb2NHclpG8PLS8Y9lOuSm9jt37XL5f5vTmJJX6FUrZdE3n8/8eP
4Rchcgql9EpwGxui0sCrDFs3zdJ5ZBVbz0HtsBGNitazUYvYOhpO5Thhbh0Q0UNnYR7pUesNSEQ8
keCKW+qoaHTR3Dm4eRTy/yaD36FkQO3qdGA72SDwPUTOu22hpa2Ox/MvEdWPBuBf9KUA6dJSLZAp
C9mTZteYOdqVVSwhaTBGkl3N6OX+VJiiPe/FmQ1E/cWETyvzTKDewM61+HChY/SiG0LoSbp70C7m
8Xu5pRnKeKCnOKlebzmIL6wObyyf/NpVYWj0qjvIlGeYYSvi1bNTxnRko+huR8joRbtolfyOTSDA
gda5DfUq+fOHBVWYFtJntR/m4SipFIleP5oRhfuK2lNu3d1F0pPM7t/izile5Pv6c+k/PGPpGbLU
11orQwt6BLud/W+9q58kGFsXVliOwCcRqVQTBHfcBjTEcOZGqJc+DYnksxWR+KicxU+h5RckCJsG
DRVLVUgaaYJ+PnSH9NMW6YAOQdCjfVkA0v54gcBV+0MYsa8k7LD4L9iiWmo+ZZrGIXYBaQrB5zg5
/5Kbrwyg7uEFte/gxruXtac2gj81JQCg2M0PuKXk11UyBe3mVFEotwgLDagssPXWe8ag9qHwPU8z
mYIEB7Vkie2aiYP21b7wGhAylW4kQYI4dxlX6p5pMPek+3LQQluDcJB38F7w7Yh+Iv8fQ18LrjKa
L0crqvvFAzZx1tWbYYZ3on7xt5ojBgAirO2kL8S3W6ZybSYfQjm1atDuZ3+uk43omj+jzTJu25HY
alcEZI+wOsRHpKuPoKujXunMk8Evj2GX8JMEG73B6gNWuEX5qQxG4Hd+1n0upKX8SjibQ+N+tDAm
xKx66nrbKplffABEgmD3QwfO71MFX9VryfSN0VdX52Zl2pFvsoloQC0gXqBIVdgCfHHZGlBfOlJJ
RLuV69XXiOoxNZgm5AZcPPwNLocC3flaTt8UOAALSxCcbASOYpGvrMfCVDQi/r9wIFyfOlgatyQ9
+cq4d1+W7nuA5o4y0MfN2Ha/NHLKNY4I5XrLhFXmgX+e3VRtpQ1aLaygGYNFPZB8KTK7w45OSQ5e
k5V9rL5BShYNt6FMHEAdLYI7ZA/PNcQMZaHNVNug45jpbKschbB+V5zKFNe9xm9q5Hb86ktDd2ql
4wgt8u8GEUprWVMCBh+DWlZF1VZKwbMvTFzVmrNHmj6Yc5soIR9gGQOAb+k9YCorFffTrq9R+5gJ
ucFjtqRi7+AEOHgPeXF3y73s9UTT9+D+XKKVQA9ADtlGY9fnk52WYzu3AnujNtjehJgqKcyEHUxv
PV/prnmPTnkoLbnREpSMsNoP7ARr4UG1UUdk+sVZrs8LODmcDFAvr1D12lWVK+wrfY2TS4tyiMe4
Qqw1Do6P2TcEooE2rMW/JDLJEdnfI7cYxovO2H+FzsfdpvdxJQqEZXRK2N7RxxTWF0i6NiErs9k5
hyTCSJTWuUKA/Y7QSAjxMzhd4XCQm3AvWck6fSm7Qu4Ts3zLdolegomAYwp83y2iiVimsKTkZbHD
9qixh0mIjR4231uW/mY2RCX/bJOWs4WgtcgJ2S0A+Cwb1wgmBE3SEyJaGrUWmeimIIwTrFxsk9e6
EX0cjD1ouvW5TF1zxQnhDA5puOEOXBkE01LVH/pROESvEandW8LGhBqeEtHYwFos6Sfc7bH8d20V
3FRmNn4YbAjHlP/gU4IQw3/9jIwASAdL5ggLwl7Js0XrJ9F+PGOUMYuoWdZL8ht9ElUrgAcFsj4u
nOtfE4M5GdJLOxLLjvXQoWq0mD1r3FeA3MYO3aCmF+YB+Bb7OwpqI1EM9T6L5N+wZMoARwEqZXYO
ZoJ0dlp/QZCf/x9GDI8mcOCqP79zCW6edNbZEnBFx0MS8uBAltS3B2eXB+/n0EHMZKRwO8u927L8
z6WNUhYymOdD3BjYOvkTfhcCWnkw/idFIZCLvNCIGOzfRKTRfmbX8fHRcOlqPf84AUQNy7pL61oE
F66JPyLRYTRfVkXLFGjJahg43aRrsOn1WP1kpAvEgMXlpdKToZNovKOURjggrRQsoJD0rP1jmGUA
kaXwW17vG4wY8QcBAuSHhA/GYgoIK0WG/E8lGde6bJMCk/5J8uXLtqN4XV24btvxE2vE63jY1vHp
bo3jdHKmdJjF3zDuJ00408F24TuEzR18O57YG+jo7Y6CioGGM2eCmysX0Yqy4DLJIAfGXfqL4Ccl
PWITAmaHtSsMD59aMn1lpo1/Iu2e6+Xv0r2n8P9sqKQbZGKSBah3Ftm7ZoTldSAuxSNJ4lIZoy2q
gWCiR3fx/M09GiekaEdrR6Hf6xaMKP6cbGh5hxbtVTMBW60EMRTFRoEj5zY6OuB/xiEqbI+1K79Z
D2SAKQZYKX/9gF8qMOb9HtXXOc6JDPBr9HlE2p1Re7kisl3rJKpzhDEsFGCmO7eK3Hyph6b8aWZx
DRAhTQM7jUpCkzI56ObyNcx9w00OxQrXV85SizO4jZXLsIPq2doEZnAJoiED75fsP/F/sAwRlUtb
kwkNdTpdjNJBsL3qgmVh9Exc+tN44fteXprgmNSxwSEdqxlfebAxRTw02c+x7e1yJlFo9RJSFbHG
xAcKGjoMBz0pINDS7Hda5P/GFBE08wgtNmUdUp8k/vSoSR1pT3z1hFFujmsBxz9A5ruIq/ogzrGS
ljccU1iiD+aXBZuELLAJ+ww0uj8Myu1hERL4IR1TGHVC+gF0o+2AsKLnVAdgDumpRq8OdS8lbTdH
0ctt7+Cf30G9l9f+2H2b/ByjPXE2oUEm0znfIuabdwtclnlOoBakbwgyRxT7s/tCWC5jOetJFuig
svUR0LVtx1EqcdGEpOpdTRDAhdjqRAoJka1E7fUHaiUCn2nMDiPLaVccijnqlU8R0/R17T8/liKs
kbJR+2mCWJCswY+Dgx0D5vtDQC0aHSw6UioGz6WJNQpWojl5HdCN+8p4t05OM6R4ON15Swg5ycBo
u3+Ux2hznNlhRLqtHGvwN5l3LmuAOkPj4lFnOtb0q0OVTyIup1LXuX59RkFdm/dHzv/C0KMalKUn
Pl08/srSfl2TYNpuZoFkmS/Sd+ZBULH8iPvX7DsKG8QJ5slDoB0vdOFCU9eo4dz9lVaVfcBxsrA1
YFBqtxRHupvftyAB2la2Tn5IK29lt/3S2XjQWMIjEgsKbV1eJwSczQn9122UNt/AbXormX79y+2t
euqCh82w5ReOn7xupKOMXX9cVWWKwF57Vf5m60HBkirbL+xQ39qYNPCoGa3Xk71Oiy8KegdwYVLt
gsc5JUnC2bFN+sPuhls/O6rxx8OumnMBwf7FMXpzYQ26AdtCSGP82RL8gtEfImepx0hqF3/ld843
ocm9RlUGjJYmX2CeXBmMseaLzVkneNFHzVNBxNdATQxvFI7oyv4OCC44oEGw5MJQCJl++dEp0QJi
PKko9gSM3uqftseAe/v9YPK9gWdOFoC52Q7Yf/zz+uhpFhMSSvjEgkYfrGy1h4gEs8cI4LutKGKd
Pvg80rF51dGK/Bh2k/tiX1CaneWfIRJJv3nNBFqjyMQW9dnoD2fIna28WHU9visa5/LEFeyog8iW
sPWgdZ3DRp6T0Kt7qXuJvX40SZpHSLvvperTBWazpsJlOMjqMx3rIu3N0Gg6ZUDLJexK5QtP2dys
bgPvnUerCJ5Yhiwq8Pwa5262nOUPYxyDCvCfNCQUn+Ttf6tCWWjdetzgDRlmFJYzE6B8aorZ7rJz
x/smlAGELbx/tJX+HljZdOJqWPWzAYvnS+waheDxZ1ALvxk0kx2QKgxbQzSFZ23PQSo5iXtkK+mb
qo7Ii0sdNofkgGb5dehCtigdrwRObzpfci5FJZQ6NJTpalYxdWDYIJKSg4XS9KGQ6svEfIbUGQIj
z89SXMpImEsKjMZkYPjbZx1vgnbmZfCZy9koI0e1mX8NYpC6WNzdCRg8S8lBMEU5Pv1l2aeMxOY2
VXFdBGSJiB88aNrpYKDQcl1Lbe/yXGNx9oHfCLFTN1wmCU6RSI149z7YxVTy0vFSEKyLfQrrAEl4
uft2Y1vqgQ1akg/LBgVIc/l94fwwdFkIILT220N8njv0Xv6pHM4pnRn9rhe7s1z0UgM4DVD9golz
Xw2HtASx/3/KfnT+PQILaUcj3x+1Vhfu4/w5jteWr3QekhCvytvYm7UNLW8kXgZu6f3t3IJDidV4
O0Lj62YbA8d3yzWOxyA9rKQOQGMbhysp6rX7+M1shfRzN0kH0qPUqD/yLnGmHLW6xjwuGc/e3uw+
gDaGCDb32pfTYcJTayPOVzy+wtqDqKvEd8rj1ZjDVtklgVMBm4D1EYdhpFSUebCcCAWGY6LGKU5k
HDauCKtZIOuo1afZf2ju+kW0UAIoXxvbIi5FvpYVCvpQug2p85NRaSkrt+nUdLmoX6BrHwap2Qkx
i5Vaa7JaA+E0mU7hKyEk89pO8ZnMgBSeBPZELC8IT4tKa3aQtsH1Lga6Huaq9sWvOWcJCg9HP8pq
mZKjX4LSqFsIKEgEQAkOX8YscXt4tcVSOuri3+/4mSvNOZgQI1TnaoLVNJzVOwB6gnS0Kf2BEQOm
iWhc4cMKz5yejO5Sf9/9POdYPIGsd7BXu1BlhwTJbIIYFH+lSxsTUlEcCrlx7eRGzWzNOoctFSE5
lP8ciuIMMZnIx8EUGRdlMy7yV/vEtGZ2ZWNyJCgeXn15l6YPBV8O7P5KnO/mnRdRZBkabq9rE0Tv
YjgZJWJW8HQMGpUole+MvvDQhcZFjSKRXrFnJSKp/1ZdjeHDlinYByfQQnXgcK8Nm29utYhYIb1L
swJ70DUbybeybUhbXY/ZeI2+L0cox64UmC4NCoM/EVBJkp7QVP8tvw3E3xB6H/Oa0ud6m2O180/n
zJIS3CgHSe7QEhN8g0CDuIxd2at7evjt6/gGtO/7uqUAm0ox2FPQQCB1tOQWPwjDain7GAd2snUh
ds7Vwk9jXcJP1x51ZLYIpw4ZM0/RuTc7P4hiNM6Q8WBKCf59u++yiAug5nGZGJ00Trfy/YApZx4X
s1kHC8Bk0gvREkor5/MRt1+w2f2kBj5BQLyEWE6fkwh+qyyH+bk0C7taQFoec9lcxc4fGn9AAXxt
ie+eJ+TpZAYDJJUuDMl4w9UuomAXJL8pOdK9BvPGZxc/sngAEWEkI2FwhUdTdanwhL1jIBP+QX1i
m7DywEXrd9Go5aln9QRxH7kAtZUG7ksJ11jjZ0O6+DZfVEpE3nGnQXrq1EpWZz7UuwMQS8YLuqp6
s9u3apeHMVZmy1OUAdE6nV0VY95VhfiLmAM56ey4RCrMuOFYF234EWE+03M+ru5vsqSThVjvCcmN
sbMuPwi31prkqWG4LW8M0HTKS3JkbjFnnJ7kQtoW8nE2tZnXKMfZFX36dGjeEM4TPjLd4F0ndDNH
tgrVaTJDA9+MY6bamLvpNYlQ54MjIYHt0HTQnJPj92oHRdxU/moyiaAB+3R77JuGCK/IldniGg7C
AAhUrZjhcSiaHZCSf8Q+Qcmr8Df4t/4I5PfHl0GRGIgxqKOJv5cttPCgy0jJ3ZbKu8LpXrTzQli3
YXcmu43kYVJWA+tE4xV/X4J1s4ga7R1YmupR/1js2p/ENWbLGDf50k91CFVfUE2jfl356u6uxLLf
08U88DK6uMyxKW5J8Q1DZdH6L1mT0Ko0ecHWomo+nZEIxTyxuV/Uke/dUqk5+oIi765WVjnPPM8A
Gs5xrbQV5UY3jb0eKxvxb0cgGTJ6eFTj+OID4oKw9FnXeOSXU0vRXQtHlPGer7mJd144/UxMLqeu
gOh9+CW9utdfMvBLZbaHjz/NBEg+bg9ptgvjsD3NIXAjR9BTg5yGozbdsOJXWnyRDBUAwnal7dlm
mETk/qUedxO+zV0qUcDKiGtqEoaBWlLTU8GifLGvaolFLzlkDP1FKGhIGG9IhQOT8dTywgUye0eY
fgcufoYEp8wGtgl6mfI63I2+RhU+h5t9i/se8WNzlnzrRk4w/yAPeJALbhSymVqKgFxaLjZOiCFi
z84sdqVgVE+1oyZ6+3Edlc7uFYVKTHhFnupzEMbSlb0wZt7GCYIRIpsoKB5qFngJXvK6xb4lTOeh
BsY7or+9fJesjqs46tO2WdPq2jzOIu73KQ+hB5k1lVZuLEO91dEv8I6FTWjiMfHbufOX+vlaXT27
V6lzjoMCbvLK2lLbixTZ8qDe21ZYnbdmD/x07UyePiHqOfk0R5t9pFgJubfPblNRwK3sT0eEmNiV
iipo7eHzvz+i40qFmtu2DBwZ3f0i4XzGZFHc2QPj2n9Z97YMjhPZvRh+vPraGGreegAuCa+jcYfC
kFyB70JnIU8qBuxHKdHyCZc2Yzi/5WwgqYo/SsfTygoqXLBdVWS5mPLxvl8NJ8ItraQ331+mAsOU
UJShgVKpSbCl3CFVf/d+ejzdRIBfmD2KJgvBmVmIKL2atcGqsZ97B/L24MzqISDgh1VRChfx8lZP
zTpshOUfe3k8B/2013fCGxMwnrXnC6P32Uyip95Bzv7SIcblDskk1oGf3tO0J9icclR4JC+DtSa5
xM6g080uAC66+4ff3YAOcdeZyAW888T4vagnFwPYrWcrF6tPPMJt3z5mqGemcQIzF05MRE4SNrDn
99HgDyQpNicH1DWKBGZ7hBM+Gb9AE4khi5I92CewugOkaDKut/ug1qgsXCpc8pRg5N8exLlUZ2XP
lgX7RT7sKQLMph5TLA81oL2933LbatWPmiadLpMaONLpNoWBR+fcTzDTyAokAeV+e5faI1aIxoE7
xrp9UWsMh2p0m6tia3Z57ta4FbwTdCeBecObuRkNWqu7WXo6LHBSZaLIcA9byzmmthJdCGidnbqS
XLTrvki+q2bsjQIOZa2cx2kvb0/JMZdLoqpxG8grDoc1XtPCoUtopy01It6eppzlwxHWz0YefL4U
nAmoKyTkVbnC1pVq74Zv8JNSFE+a8d7GItZSx7w+ozCPLdO3aMmR2H2j9mshecAJ4P4XAsOMHrDa
aLLEJGCAZc6OddW5eodFH8KUKaUgi2KigCrQ7QjXrzlS5NDkfZG0hU8wun5rgzLGikUWYADbpUAb
SDFzSCizxEmIyAElPrS+gHSJDAC8b4p8NQVwYA44I5U0urbgsxRzezQHddEm7+vazT7yMv2UdKJV
RtywJG1Z6nJxGqwn5ebQgBpK0RXl45kECdYWNo/ILFN+5y3O2Kn7f+EozsaPWGaWgkBoS0UftxSm
v6T/MfLuv+QtXrGV1Xz90V4mMJlAgyuWPLF/ulsSN5QGqgkyA0wd053tBdESdFotNeD/T39cd2aT
PzIlKd0slpYHlJBMdoDbP5/TpW1Can7KN9hresbrOu4hPHs1gMYu7zsWNE7KaZcJ2QvqkgAu+Obc
CRxTWxSQwneo7n2dy5WqfZfF0VME5c32ZU4xS8viYV71FSQaryjAewBeVC+TZ6fXcgiUKTdO6nnT
7vgr3YEPhurAm/+QFYfTodEGiwiR7ouoObzYzYhCmt+wHK485PpqJmjWHif88ZCDlaIx+m/MXdmU
z949q9h97ZOyQ/ZHPoa4YwDzi40dtCsJi2PH4fmltdi/PKwWdVKPn9p93oYi8fi3P/Dm+ZJAbLez
lNlBPIpoe3yfNxscKIr++Rw1dotaYHpCKC4uGVrPiiU8Uk3VQsTemHzKzRdiEPP13Ycqsd2bU/YP
bSoIKSkxK5SKGDj2L3Jeo1LNzJ6zld8Fkh5mXA7NeBxHbXM2qPs6K0c4pKXmvdcxUnuiWAy3l0ZW
kdu+wwFRW8vM+nTozw1wMdSvloXmU6FDrTAZhUv1bQooFKaHiCMVaXDmY0SKuTp32AyLkeWoYSTw
1uqP24HVxZGgbBYx2A0VxP2/gcX8eH22T8363mH3QguSxQFU+g3hzwIFfWNKYgkzEUbtH5QUVLfu
k8RYr2hM8/6qFpXlxoqWlGQLKE4QD55O8DOoq16iqUfUiePwgCGlgZhxJLMfyP6+G89CTp7XwOI4
Q6xzA4Oh2GGXGhFnDs8gBk0nOKF9g+LdFwM1zrEG7T9NFTM2XM53IG0zsMcBlV9Vdg+UZ5uY/hiv
2vt22QCI1WClCvWvY/rFhTRuXglWIN0L4TX6fB0rs1aJ2DcxUVDKWibIFhmXacWjZGrMnjTZ0F+7
HRwv0woFhYPRri8Q7rCMUHo9x/a4XsMP8BDcJXzC/dzlWpu/pGEhnAIo7M4kPx/qvhDOkLcluD6h
kSNqIRh0EufykqbsL/xLcTwjy33CJ+NADWkruGnkfunaTyQK2Mb0tXpMKiJ3lZ3fIaDkPeeCWAJ9
yKe/y2MKLMkg1MNanJ3XppkYaJMrxjRM98GCcBQKvjtAO7mxYGBndp5Ud+da6Y+5VcI6dZRzB09u
H6h8ObYLpDqjHsTbsmG9LPmu1LHoIh9XEMw+ohrtDvnXB/212Gu6tdlFLDJ6O2gg3e6LVIqmIuJb
vL8Lkzgs1T4BIQsnB3f/7FZUlWkDhDtdAl9GSWw+8voOAoVb5O2BechxBOiKZzcOkqcMjnO6SpGo
bveVIxj1Zrbt71+7MEE/RN53Hucqq6CgeXb7VfS3AC3c8lCREPIH7DtogiyHn86rWAIoWTwBkZNn
OTyCi4imecoFXqN19z/oHpG6xvaCmT+ljl1KRSja4F9d1pD1YQY/KbqPQif6FLISHF0YDnmf/de0
n3aOtVsfbpGbhIfhODUySr4KzMGHCj4PqbAJz3Ax0x0SSOCSmmLPDbWfEASaqpQ48raJvqjdz06G
yuubSRHW21C0XSXmnTqBJw7guwFxB98WonluHb5MweQeM9mzOX1oQ2Jw5F0x/j5qKg8g4DMEgKdF
JkxX/29+yOdDRAlQr9/KqnEkGZELqKVxGPuCWmMAC1v0dSoCr+rEE5q9j8q/1/oC4tv4MZIOUElP
g/12DMV/fV+3SraQKj8i1TA5jx7cddglVVJJbTUskWOwV1h9x5q78xk+GwKBygl9VvtE7NQoAAEM
PKLFDrYR3x8U64um8RUguO8jWiCZGEj5RmXKTx/UAFoDIm77xIhipvee+dd77bSH1tGkgUfq1s1u
sZoCzfFYb5all7WjdMt6xD3bHmv7JRc1qvZ14Y+ExCXEFc94943S4zv9FMvkLtto/4VVQuQd9ku7
6UlnTsmYEnIuG3Wtt/8zeKaAnEnr8wT7lkiu6hZLRksCEJhJRe9X1+S6WdrsII/U4CWXyTpcjBHh
O8McpZVEY/K2VLFaCCHVwwg3hhyRUqJfR7VVtARL55Q3PuXOztzQCA7Q2P1qWsKGq/HgC55m0ds2
Y5hEy6xzsDjnR4P0VSdtuv2Yas4JhFehVmh4ciGs9KQV035oJmWIB5Oji5KKvRt3fqJ+s9NM2WX5
oOktS7E73CxQxvuX53u1veZTPT8dSIgrcdJtBD8QzRfbfmwocid7rZcph7xHdk7rf6Obdm4dJuE2
zofDyz0XvI+KnXzf/eFYfc/cXb4lLveN8baB+g9fpIJDyjHekZHPl+S5b6xruZMuw20oY437EmO2
kRe3qL+VxvcYgkQL1LnOiEs0fRovAfQoGycMdiRpdQcybdygrTMPHTWzc2eC8cfvB/x9ObKWv2tL
nEdf5uGc0SDTf21/Dn9HwqPbXl0f76x3F0QawDM223kreYCa6+QaqO6ZrHXeqjkuKkvZqGMKb4Xb
j8yKx2wTSlh+VjphZW/lZp3AAkYe3kMwMy3e2gDgDr8Wtid+iSKRaYNVuZPLPpAvH77aa5wmkai0
37hshtBXcPg1Fhjlu1jhXWqd3K0CVSLvtTDKLnxWRukN+F/P6d2JRpQdWBOEALTtXMkozyrPiC+E
Fk+lrJiTfWgycTwFbqM8XrI1zMhGulMDvsGDcvIkmzPSQfDSp+TvZiMNAF2yn62NSHduX1a6jPLa
DQAZqkKYyNCFk0tqie/MgBJaGOuoyb/j+k/V1fEiofNQ+LWGwTpnVA5FMhxZW+T9mSzq8o4emxIO
dEfvcUMEiTkIQTcLiTn01nqW5SCMjbqEQj/Arm4swR56kbbll4krKWORuTQi8kftZX965CuA1KPf
6ITaEec+VBgeA/pZwxGy6xMUumKn49HQOZ1EzMlZ5jtXi9dfaWqxzc+Soi7ntAIjO/ZPI9ic3+6T
nK7BLftGAyBwgZaxL6I+QlNWrdizn2u9JVEbJ51efCct+CjFQmAsN0N3XWGi1fBliirhECx3fHPs
7gfBmG2TFgNoaB4UdRHlbMxqPpEwdjZigS1ndM2Mk4LAPTC3L/llRIrGId8VD2VsdV9XJB8tSnQM
eiSa7KWU2t06/cZE4Fnn5p7NkVzDVp4V4D45s1WpXzLvFFW1+5bcyUqVIIwFofkvUdS4WbZW2Uqd
ziEYmIFp0cXgy5VcCzGQks/ItdsPN3c00J4MTik4N+ZkXjl5nv5/vVcr+PHq9t5+mbB+vSIP5dZI
Z8f8OQi4gAZL6U6oZZ2PXhkMhWaeIvUYWs4z2GZnBFWNCEvrVa/BvaH9pEtUzA5CQ1CtBt55lh31
dTJO4wGs8tTVXh4nX68Og1su1QCc5n3EF0njOepIdlP/yOqp1Ez9UJZlxxSQivCb8slUgKOTTrw2
uhm3/TKwnpARCKXNAM1TONpG+qaaVqRCYO7oHpHpsOw+hcXSFYRYPENMBMIYx/pfCXIQKxp+UPwl
AXPC57QsNmd8v8TEflZFGH98dhkr/1T8eLe55/xpRWT95djrLPCJLiLYGtMxX7f400WJHpJj/cqq
4rxDo39dbnBnS7+QCOnMLqlkDlU5eiymB0LSJ4UpguA62xXu/ZbjU1Sid1r/7Hvwc8QphUTc5CWa
IepX9b5yMaWaiNSNdMgo+re9ook/FE91f3LnFj9YXQeYIyVWbpR0HzBrQdhmgx2/2qarPfjIN1L4
YEUiAJdtw/XERW3NlLBd9Rt6YdBKyAFEuMjzCa48Anvad0Qah9Re5elGQ7LtPGHcg0Y/32SdCW3L
/syK9XlF95zwHbxzK9WYYIusT3kzb/hQ37V3z4YOreNi5oU9A/1W7lt/r9Tqd9pKqOpJ+5QRsnDa
Tpd51MVYgnf/AWnQdyyx/ogJZLNCi3098MB1UKhodjRsokdM7HRgjMIQoE/GqvmAWPR9km6opnif
OZcsBlFCyF1udVebXgY8QGuPAor9le6DJuhnwiGVuOvmXef2j+NZquSHZKOleWKlNnWWKNMsfzJU
5ity044lMORwSKy6UAKL7lHN10j5tcqztuMzOapaBGglN3us4irhaVW2MjHhxF7vEZLeBoSpCZbV
J802UhrbuanaT5LCcaxyUiSaMqVZV4wlgrvD9yiifgXGu2J3bGM6+bxkH7sf3eJZa8l4q9SUPCDl
hoN5DRH0aO8qjyZBUqvnWbA96OyKs8xkh0WXN93TGDQdxZ9efZ5lt76sQvLDjRzYLFh1XtFOnRNZ
lW7FDNk1RPmPlNTndknIVzFTdMtdB5kavJI+ocvIH/apiE47f/gY9NWzkHv3SsyhAQxR2f1PgdBH
qjLF1/EfvHXCJs+Yc6wNi/q1jLZ79vX+wSuKeL+FpLRDS5rfwwSH2a7kvEAjUBRT+4aYrUK5DdjK
5zj1VNZe8uOPzDzuhk1DGtFEaidlUSck/soJQQHISBdSH/8VYr0/bhi1qocNGqi1AOx6G3CeUvxr
zoNGixMB177KnNp6FTv5lUvmsuPVZdIjWCTudfk/ufxS6zYWEtifXXW9/ybxKmA13T6yWxI/ib2z
h3gQqt/tV2bbb0m6PTzk+G9j/f8MQTi8wqj3F2xfoRaH3udLIk8ZiaCpbkwluJ6skPE3LIQIWaY3
ugmE/BOKcNVxdO1GIwxQmBTS+pFMK8H2ZSkBPblft5SvGUP0GZqlyYXs46ekAhbO4NiMFWOvp4ln
cyOB6EwYNbRcXO91TLy8jTCd5Rrizkm3G4leoyQ3i/pGVupo8408Q0vkG4xiK8XPJWQg1mRcRwsl
sUu7yQce6r5P/a8UFB0R5WjrykHOw6rDQTGLBucTd0ynoAgmGDWcSJCKSANITd53rgPG3jKZxPzY
WkW+i85Fu288s1FQbiBBCifujHZ7A4ItYJC5/OV3CfAJ9Xnh2JP9nDNzd/Pf0eF9izLXS1WGpIgT
nkWXb2OdnEaWkgmKPCFCaR8qWkjnXNfWKudeTXVd3sbIZTq17c5HpN9w4PQ7Fz35Z7XBFtQl0rSJ
/OOP2MfadLlWvXbMIwGOpgy00pnGpT8REaGPwhCHADWqZ37igAFwFn0o+5qSWZsUJoINqM1K6HYC
OKpkNAhOJyi/3tnZ0PITvF/m5VOIM2KtFhXM1icSPJekeqiww2kgVBIpeDTlhBQRDgddLx9frTbm
SIl3gsW/ZoyI/RyFcGosvl76JL/RqOfQianRqeJ00RsvXuQ0OV57iOApUnVma3nq6p64IPLK5T6k
Zm1zZ/NsbDleiFLYUTvpfDdPUvHS37uKYtk8mfZoQPPDYcska+meIlSXpmO5odtatlKZhYJM7mXl
rxnzNLqaiICZWs7wHs6LoQjfb/LYRjgoeee7Dz8Wd4zzULSJsy7PBxbnGOOV76KMe3vPdrxh316B
NZzpypcdhinmA7SfVVxmUqQy378pim6AKp/hDCpP0GUsMO9p9Ow0p/FASVjRLYA0iMnC5XKFCVOP
qCVRcrABAABqe/kh/qVCpsBkbx5HNk1b2XhEHb7evN5toe6gIrGVy/uzIpt69xVk+QgZzIiLqaSG
imwa5WPzGVXIizaVZ8bYmvqxHUo8LGoraKkCKVinFC1UXJEvHSgTv9Bj712ySbtMAYqlTv6AILvs
LXXSZ3MYIULNUGHiiKoDuyjcfhUhQVeZbST56Lycb0NvSP3k81H64xf9io+J7ewuDEWis6xBSqu8
94BlFADj0Jp+ZKAE1tQvzRfwOv3f2yTrVtInyI7ZHkz5XkR/wYJmvy11+P1r3Q6kmCqGckGbeEdJ
AbxE2OujZABLpNqmh1e1Faf8NRKFd/FW9nHkhjcMGIuDogsyyfN+rbpY7bpGK3MC9ddz+fdGP9f4
jA30CRVeutePbl6NW2btDobwvHL6WRWHsfJhP6Z2BIbCPc3tdEP3a1MURM+OoeSxNCWIyqFA69WW
MNFNuvQu0WgHopmrHwuTxZm/YXhcRcGhlwGPUJ+BMDYLr/4ZgAueUlNCHwrh88z1Ud6oBrxldhOz
D2l/qmmuxRXqLQ6z8t14fX+1OhFiiC6A0K9UWx7IsbBiLBVSwn99rOXUbLoDNu4vagdeqQYvvwFF
JOCwPs5oY4UAdTInDEptD12AYqiZeP4XzJTk+eYOeQt462U+eNSaN3lc0iERAkBtb2emLwoLWqah
PHEM+umLkOdM3PZsHPhgQDWbQsS4v1jK9FqSJiD3Eh35ROI91W7bRB/1dnUQo1WXOAOcfGhQ6ErC
ye8WON8AAsWa7mID6voh8ZrLcZ8oWqPpVKDYCvrG4XkRfZ+RD+j7tuxZC5O/0nq5uXaeGjUDUU25
yzG5Y3yIUWIvddSPuhxObAxKiPdkMSKcjNptLbSUx7GdWbqc0FN/LlnC4+gf66ep19PBc5Cw90eq
jFHpJ/hk9pShk1N5nUyoMYy4cRaotnQWaReSIF5EUIZ7/Ki17+pDvgVrmlAXpE7cvpVs33An3RTK
h5OzIQbHw2gA3KgFgGbJp5fO8vFKRSxYenAkoir0alHEtK2OPSkxPF+xV05WK+V7GwkU8DOrxq8q
ZYwA13qN/D2T8F7nC5UWFGzQscBMKRTN0wxu3AOK5HHMp3ODddMGzFOdpfq8cjhR2I2ME0hPXjHO
Q3xnfyGvBHzjvouCRC5DulwveJjvkZWuEa+j46zrL5SbUa1FelX1zqDsSh/TRy2K63AfV9vCMhSK
iUFlbBobDF91m0MypWpC2VRwA+JTKFtxECPl3f68iPFqPp3Jx5kCz6EZmyOtGoKHfDRNjNn3bt1K
WjwSFLeWXYqHRT4irIspeVhAxJBvlrUkBH+bCZrj3nOmDOqtupqQ7jHxly8QqW23ClgyCKHP7O6x
KGvM3agb8D2SW9R61QKn3XFAlGty8MS6J3vDyg/HasnboEVN+AvgyCp7UXS+Pjf0eDHL0G0nUbuz
9r/yHJulWOSlSMr7ihVtvquXS+/oA6YG/ZCBf2pZIJySnx8u15rk329ZEOJ2KR+dDo/UoW++Dpdz
B9BTuy5tlNCHAhrXfJaQxYLhwhkaiBtnZ4o9QnzhLUQqMC8oO96dSldXFBT2sn8dnwrBNKSSSutJ
8+pvyoTjDhu5hA5mfH6yy7/mw6ALYg44Q3MQz3tRv4wA5fmlC9Xonrwr2Raj3/ZQTyQO1444LjaL
QxzyX9L319I7CLWungEPYKuHXia4Psa8uMYP2uc1Mgx93FsuWlUlQWZkziI6NEmodbgm8+w+/N8q
1Re7++SSZ+7xGeili0+YE/nmwNmoBVV5hDCwwpkjwBVaLszpkDk199gnwPP4mPKI1Px2f6QMBtDZ
KQN1NZDbqRyAIKlIfaa6spAJUv90HXlZKdsf1ugyIlVVBsi/nRFY3VUpGXyMn6PYv26YJ2qRhpjL
vH3wE81KiqtBEOzqVPuo7/5kj03b40GT+12qb5KgHQvL12SuJDh/VCYPtDI2ffpaXAhGKvcfXIjF
djcVRnxFSC5fDFnvcRfzq4njANq8FJGI2GXSVYLrxwU2PxQxMQaEcioGJLFDpn+/PFTuTjrJoSNv
6chjyb2pMCpMmio0XLceMpyPe5JS7L2SYscjhcu3+lwRKkqpzuc+Soj6swz31dqt1JduZMn/fnBC
7Bj8DP1omXc4q6dBtDkMf6ScRyu7uqRoIw6WiiIFsAwHyEOx7/RV3qYs05m7rwUXeCQr4jjhncE7
8etLK6RjBlJIMIKyf46kF5DubPdu2Ao41L3URAprWGpSeGTnzcGRBXU1dEHLlikHGOcgurWSoLlO
gDZY7K2/P+tyTJSS1psq2+ckbuuyjqVL2HAaYFNCIptgisAMroY6opAXYIKXN5hAOypNdby4sDxE
OTi2oXrl+OUwG971Dl+7okisUJKEn/nmieTxVmWuDwHz1W6+HD205UFoNWJ/4vWT6b1gBspHSQCh
zNorPT5wIuyyOkOjPHalYZJA3h2knvPwsCqX91Z42HLE8pKFyapuSjIXc2j7HudsZ2eEtv4lM++p
jUvTNkC9O1uLiGo1ljWjTPmnvf5g7Ho8T5rgdjtT8kpykgTV9jgK55zmHs9T/AlU0I3cy/Vc+4BD
zNAf8fvxwKWsmnOua1YTcSw6t5w1MDB85XEBqMfBksDrDYEziqK3Z3xbhlHprx3OZZP9Ck+CG5Th
9DsMyOqiu4rkS4+nH5UF6+BL2EoNoYN9M52mVZuGfC8qnQMj1jLylO/KZpdOWmynH6ikpnJIqAhf
1w1B8rYXcLNCrLpK+bK6MbpozPTns0fopclfWTCRhBqnP8Djg85AOwsY8oLRA6TSwFXic6Rjio3u
9KYsLlpFdCtqfdNwtJwNs/CdFxsRS9+V42ypc4JYZNrnVpMBLbROFEMEn+jd+ddJrNUUTevjId1T
xmsFtuZ3GOjdF52BZ+ACdUAkWXrTKBMN8T4HwUrxD118Y6/R9TjwF75oK1N4tocbpzf+cG6B/kqQ
JH8RmZO8VovbOuWj8x/QMC9xFv9CRDl3BMhYX2/yeobZ3g78zSO55A3ObonJgVq+q6iDbP4s0dkC
xelrY2fXExvYasd7rOspRIbOHWL8TWD+NYdks62Ps88PqccY6n02wJhrRnLlXfgv0lxcqgP+e25G
TFD6FI2/dhkyLf1f7a/4fC12RxLV0aNJqMerX5vOiZdtMoyTB11kfvg7l6BLO9w/ulSB2fmbswvd
BxxBuf0q29h+GKFufL5VIwmIIVzSfGwhlfCOtEFf+SEvD/hEgiOTq5IErDhN50DnvFawBBrzyiZU
RqFH5jniyVnreaB8+3m9262tbSspxJwIJXiRfks9v7ponYXCXNciARgY31UlmUT+TNpajZCbsFLq
gQ61GwZ+HeRGpasHX9dUn32NcxTQCVWALduFwzulf5peFRpbAQJIYIChNNNjY3yYyv3BsfmQFMOE
k6nSa5+JGFrVRimagrZSGBozegA8UdCSjMSdyX7j62c/Tzka/d37V9+O8RiF8Z1fNXzQV4W0C42P
gipq1fWMGwIkP/RLqv2uzlCvQ8cJ0GZH55lMDh8OudG31Y1Y/LPC+u8ZOhSkH/98XvX9a33uWjAJ
Z5pm3OOBLSyi6ccE2MJk+FHPMysf2e43drUD8QL+XHVqLrS8z5TxpltFMajP0VT4L7ambzpYEhC7
TXtzBK/stxZOTPl6T2dGX6fbd4/WxfxGgnIWzd3qSM0sOTH3XEP3pq5lFsZZa+6vf6AKnBlavk2S
iGLovbE9bE0Ma2igQXO3WM0bnXlFVAQJa+WfpTAH8mTeBjKEN8XlNJF6XubPL9yQoegzlvoqrQ/M
eC89oR5GiWMD+NHUbNzpv1cVtXi9lv+FvTr+9K4FTJ7mB0qwxEVF8s3At2LMlBffuNlhIzZwhIsr
rp70cG2K8e0T4ZmAk+kRWK3lpAjIrWpyXbcaGFunk4vd4392US92XYM63i7ec6v02d4KttSoB5Jx
s1RnsUlL1fPDtZM0OZR1ekNOv3iXf9mNbNCQaTg+Dsrt1ZGc3K9kZXukAQMx1C9TLcSZZnnz3trG
fkdqyjXbW4gdGc+A1T1ezeOgvqqCYliiEjMzZc5TqM25AOjVAbbhWxZeKEdCyFMROP6H4Pca7UqP
AXRObyab5dVc5Ie+VE3NkihG31miBKJsdZGHOKg4hCGiHJlCnUMjKC1p9DsXpc2Jx4/PU0h6+lfZ
/46RXhlnVMoBpS4yuLnxgQQVPf1ypppLpmbE6Wm2mtTIiRBm/RfCxZTPS2op1zsPa7n3qdHhtVXE
EO+oeivRgI1t2HRSJEOiWSunbbpUuXjzz+yMMXpWWtTqU61xkqr27/2HoDBfx+JEX6od3uA901EK
K5NqwSDnrb8Llqgbbs4SLeRK0+7T/8biQ0VRu6EcOZFCpkmwB2XwmaODgglD1ODIBb5zwbyGsA24
27cZk+Mo1qNDdx9aNYsplOOZt1tN1a65hrX4X21p/RVeDyMc3wCEA/ncyN8DOlOXqifeiNTFWwfK
tc3TvZwpCUycuKEzdnFeozeKl2ATenR6IYs8H/1nWDgiPzAwrgNYDuvTmwj6fJpyU6A8aXyiF6Sa
4fuPZ65MxxqsodefwdpvUHQCd++dQ/wE/3jEIFv9pJIGal1xpvsD2pgiOeoMkxVFa1RDFlsBerjQ
Ppgn/zzQokS1k4/DQ8lhMMtaCbqe/ze+PzoPfPmB81oKSU2NMBAkCBUw3oti2NbvYYiEn7sm4eby
operG6Q1OEueKL6o391L0MWq3u7YN1Nad75DbKml3NuK4CHOKbnqTCXnY0apmwf1Pw3Ir2aZgIpm
LJAf/1byons3W94H8l9qoa/LQLdWSAvW4cCSMYqeA6xvYrPYcHRaXkZ0lVKwwXI7K9K03sWvFtDp
K5ZE5vPfYnyraGoR9+CJDMOS+6mvtJ0N6H6fjqvC11YzabVJ92Kk2G1Co6Km6NRsxY5C8oJqknsU
HzkM4Je3R6qbK4NkR6m+oTLKUe57uR5RcodOipqoqKgKj2Z+Al2EaWZCMSjzTUMInZD3XIIvDawS
0bHrVKJMFxDqLj7WH7eNWRBL9QYBjM8ExDBy338m59Z9zzVMk0xYhlq+a41Ux3raSUlA6TEubs1K
JvSo5kvHFneVWbZViZZWSfRTr0JE943z6+SEZHsQeAaCjcT9O8dy96/A++3sDsuc6vKyMsAhB9uu
FJ9dJVqx4X6kDPrdi71oztc2YAB/zSxRrJIf0u63M3v+7NGRsIYkquxIrtF9G0Wzp06hP973uue5
44+aD0pegvC1iFeVhk2adcTb7iyQ5db9Hn5V0E1fldwpyg48FcBJze7H6HHiJu6rPWaE+Sao+MTH
e4GFSTLGAw+5CjG7rRH6jp3Q7ux/a7UP5l5xLxTmX8yX+PqNVMlOi6vqM/jaj3m/+mmx97xdtJws
iug2OuNNkHHYQR4DbqyGa9WUm/MS+sE7BUAVA7jgW+2toQPPECO0p7MKRAVGqPXnwa9soONaU142
Gkm6ZJdpL3jKlvj5+YP9EUlICWbAjtju9H7wBFsCc597X5QCy0WSSoL0BscfDrGOb/wCyhRs8zkL
12xu1aggUWILkws0gWVx66a2haOXy36uIIC9nPV3jTZWLD6/ppV0ZEo3qgOsC0alRspkrKf6pC4T
IXYMWwWuFeOavuTX7XuAV+W+Hvq9l90w3pkFUzS+zAUyQChwkPJ9Bj1J+OfzN2BYfqDmJz/6OCnX
RMBy0zyUn39ry6omkUauAc063IdRqGsHu5Kcv/5RDkPneFtcBztaSPLnjdqzczV0an3LgI0IbN+o
P8gC5zw+xjDEkxVI9Kd2iOrof2KMDmB4Q74t+fNwsn1Dn6ihh7VF+lsziTwDNDWHYFa18PObpT/V
H6QI8lGupFhk7zm33NMmqXRiSkcEccsnpnMCaf5my2aOq35L7RMpfq/bjyiDOLaz/ipahYFRkyzN
uAgDhBkN9hC7EuH3PdGbcEYfgkAhdnMjdK1fpar7/ovVsb/Wd5vwkMcFPNWfAO6n1oAfCKVPXEB0
4+tNOY5uSG+5qezA4l/KtzoMN0DoSSFbYAAgh9Lgqh8EzK1DxZXMq77G5t1Qn31G9UKbaSGSLQxN
8wdCPkA7duHVjh8F0NNGz9/yT/1MJN5UoRlyg0MZOHJ5+6bP4H+tIt303sn0sh/fkUF0dFRtG5SO
rf5LdVz8X6+eBfMnKS+oHX18Wu/sBgdGGq/vroDmGTNyArHUP9IPHP1lvLVUkQOkZdv9pUVP4nFT
UkSZW7INlqf1aepHTs/8bP5kr24Qs+izeU/4KaTild98r+oM7FpaxcWuMuZTW9dJG+XAFqGDtmA/
WBPP3wtvqGcZvEvu8XNZsGJx3oySwZIyki7roE/0vnxsbAQKxUOg0cjCI7vlTr4aYyvTCf0MLQir
VzYjMldqVM/7PH74cewbBJdsMDkeq+p/qGkJyOCTYqr5mLnAh5/UWmXqExV1nDP6vTVE5CslBjBt
wAboD578h/8k8P0nYnycQkhwObTgEEQJ4BtBkov8huPWrtUy8DPBu/GpKNDKj4VXHYvmJrh9wp49
DzpRq4K4OEFq+JTl/hl1z0LnLO8kXUtGEXLU2OszLSa5ldpH/iFAu5CyNhDSVUq+RXyqOuyzaqcX
H2RJa7YaSwAc90jXmzhvFq3P9eN/uDIyzHVo/M8AGq8F7B0ndilEhTIrjHFBAjNaUszx14lrDWFh
vZl3J1LwtmrpCrGEI8NNhrFYbTy07PvdPlwiEgge0YMSxKtYDz8UG19LyQLIME9ihnfZRMNZJ6Y+
Fd/zhB8DubIaQ2SlKJyYGw6Irryik7JH4Y7xI/POuu8ebXjGHgjuJoc44X0JnKlWkVFSypvHN276
3ORHCt1zti0O75Eq9BlN9uP0FLBIWMrVaYN5sSN4txmSVHEWUlGYb3jKNH/EvLvNXRNdkQehOKav
tzVYAimplXVkEkRw0CTnw78NiMqmCzRj4uN1tA/VHtPpI3oVn1RCES7RU510RVWGIiX7XfIqmnll
SkXz2ilAhf3HWl4ga0G/V8C0PgtmMcL7raqihVt5slcqHLgvhPltOL+SRvmv1ulB+UrH43TUOOYj
c2cCLlVu6yEFkKqkTWl6QWPYPOtCKv+Lyf3rw4dWwe/2Kz8jwlKHsvoPRCLxA8uTSBAbZ+MmMFVB
3M0gnYXzkA5spFl5RO07gntVUDy3pHSEHRAvq4EEMJzelEyffKqIwuvslPWz/YB3ia4m3QYrGKyv
h9W9eEV9wUAh2GBCNjpauwC8JYInpeC0/ZFmc7kfnVfrYfbffn4BKXaWmjVLewt2SfpeEWsGloBt
LyMLas4iezLMtq/6+G7XLJoHJrsMQ7iLa9uEsl1RBffgacVT276iVLOQkN4fRzUdU7x+LvcLSPEr
YkkmI2o4jOPm48cB5+O54OzfD7gmsq07WDE1GplBKcALeXuLMyF/E+S3uRgNIzF9n9YSOyIaryvw
H/22zCPZlkRaeqKkU+uoGoiLzkbNzNHHnsyK0ETqH6AYFYiHIxLuZQpuAcZH6mIqT+5PYV6IjOHS
NPpP+wagT3Y4LTSH/dh8JjO8LA75ILjyqWvBdRvIq3WCiQn1k91p+yMRkZaPzI4P8tetxKY4IBwn
X/IenwtUPf7Cecenp0a/aGotC9yJSni13iF6DfC/kt/qEzJIcAbUc4XsbZ4KeoB1d/hHjBsn+1dc
CS7vOgCa+pwB12Xpx3NqIGQhivkfcGkDJPrwaFR2sOCiI88X5tKX6DaW96ssSrgI45ZTAuVIg1RJ
CYdfk7RWXU4mtPyB08dFl+QVJDWjUmknNJsQy5uwPRR8ReRYfUWHjN5/PDxuDNqseNmoVp52bNnW
d86oi4lE9uWpFJCJ630JhZlx1iuyhPhrNSdjInTckroRGnGjeq2Icrrh2Sl6undGrAlA19IbQSTj
rTDXkUDkT9+066RSt7gYregwkqNYUJMN5E4icL1Xa7ixKudGZMzk+B12cJsFZryKNCp2i11l2X5+
t8mZHYJmUJL9HnWYyTrGCCHuMEER4bDmAATHzMAGgLFpmG6tg9Cxn4cZrV3+e4hJUpZNR1o+Z62m
w8e2STbb8h+NEo9X/7Fsm9cxWkzqMC9xB5457o3hzF3qLdgysg5fveb7WCGqRCEcTdR9L12dt5qq
rgpOa5F/lMMEEzsRjdHtuzC1NheeByJNVfnxwX44xPr0uzeAFZyNvBmYPJ4vjZGM7yXOvC/rTbmX
KSdkCyyzuXSVVVtf0UxguDh5VUlAoHE6EFKJU2EUugnabTk3h698ut/Pl/+BsJoM5g/3oWVbPHTV
1rjBfTRFzKrCITultypsu2w5mDPBSwSNAxDC7xtGH+De5xAmYegEz+GMjQlycPg5keH/E4sb0/w4
Xh0If2P+3EIuwBUR92GNvdhtoOsSsnJ44wXRRRZerKK1WxERenXksu9gVGMuNFykEaFNrorYFdhA
CFcnxFKcBnuArJlCPX+u/b5ZaXYHzT80IaCDOwsk2jbvgFHmdksd2jphkWTf+he1LC4ODItEGPHk
l+OkyiSlw3yATSwkMZqkuoP5FI2cy1zngYtzdZUBEn/73kv9Qh1kX/YlMJb0Ac6XIF75uis6EwoF
dBCYLfZPP3FeVo0rmAUilwXlZzw8AJy+04rodlXJRKH1IxJPDOJmq1ysAb5zWZvOwZiEFllH18cq
MKBkRTlc2hnPwGduQNisLvjCxvJb0mPAJJRDLBtl7f5PGRAmt5qOzR+2Xc4RymA220gG/MwQ5y43
NFFaSpDMKLsYXOFPfD3ZEbHwCS/NdKfp7p1Ph1LNqZzt9O6qK73O2efs2Uc+o8/XXybnH8aVbRkT
lilSkOKtNyzbglOFm1JuCmOEYsRPRo92kpPKxbKjh/lxT9GEOZkcuJdYeyXcgVHfk55EDJjgqiPu
vzn2dKZi4NFxDmQFAGzECFQPYHJTRzSLjMsJ6aCd7NpemMoP85mCKLrs+2sbRKRsmJWlf1WaEckf
o+eF7iOD71p8/E+mKYjwik1YXREV5lamLvXdxloNnorE7X97zBgVVv16ZbkpNLVkuQ77+/lKqBPN
E6E6pdyK1i0NUVTpoSkY8qELm2UqEuQEEl9dkfHFPYctKvo4Yt1Wj+eE/5wpEOE0gnUldFlb+9j7
KwceIf+pOcFR4GDXw+EdWvg3xbN9163H/x93jq1reh3GAbiDzGr3fl06PGBGOGqZhcWOYzGpQx/l
geFCUluOa8YbLQowaiDFDZYwP2Aaw8dNtjSeLGKtOZT7QK2sNJc1I9XAdhlWWtwEHqwFkNJjYKFV
RhokMWetnC5hU9rkG/z3W5t/529eutmVmbrpg1ZbsqCcCiy9lIMhkzD3CWDHukhWfcODrkcGbVFO
32aup/IylA+clBp0AX27o5R3JSIZIFcInfP7xvf+zcNtlgPqp7FadUQVmsqhsQyuUTePCRDrUZKJ
bBjR5HNF5sI6ywQTywb+wBU5493T6S0PBfnqcktyc03ZQORJLXgY47gt5jTAe014BZWDmgUFHepk
PT7OjRuJcyCER4Xx0YyWnGI+sslMD13H7+a7Cez4v0y+KJmK25CCXzlBcc3ObXQjD/P6S/Lv90Lw
4VdnVNpz/qa3sS7RkROT1vFiZnMZI88i89jJmNOHSj+bQ2QqOlZ8GzTNorCShCVWI7kZ6jq9f/zm
lchBS+LS8tbwAlUW6kT+S1RBb1niuAvEmGaf+sCFGjMvKuy9H4Un3sg+PpgdUPodZGdC16k2eBsU
luAsC1JFhgnwY94TjzEX/ZG2EFydf6l4raeF0Ey46lmwGxS472eb0bjp1NkAF0ELROeGVc8KvdB0
Egax7fw8zXCgTuO2NNkzmZ5UGqXUnsE7hTO8Hu8T8GQ1NQrOZyRKh+EB6aI+i1CKWdJTfBBMDMlK
KFxYJtgUesoDqE43U6fIAUbY5tHNOaSSnZHc2efNVVf7SBeW4nIAcfsuFpAvFPraU+OTvOCrC4Vi
WNRffJiWWvG0vySKa2muwyJq0E2P1k9RunxemauhfQIlc4K35r5zBrcSBImNddWgTtF1yBWqBLn4
QoRdbOnAPiDS4wokLI7fOjeq/R7dilIUOF1uWb+DstOHtQ+aORxydTTr7vSqZsqrjs3cJ7g9XFQO
IxhL4u08FRpTfGPDLSeO+qBh2M+12mF9rd/xNgkahMNyfNvQ882H5JlLzCMIpA6uT9CC4y0RDaZQ
D83R2FiKwTFNTOZg1LQhoFxd7NwoRLwJoMfOe2maskkZTAGaGZ3UmhLtHGggEfBNjsA3kyg1CQte
NldwqS9FuFc/CUU3G8T3CtutBwPZn/AgqnaiKvatW5yLi/r0Mi7yTHjFXgrahqlNx0cThW+LVAhB
LiD1W5Vr2cR0mVKsiEB662ceUIs4V4aLdCszoaTfTDaXRV1FwbLH24vjIKWuwc4fgpmp/tpLbJ2R
cSDtFlKKOWGftGEmAfTAYF1Vh4Hrb6zvQGvXvfMPAlCSOoUBnnTvcLquy+2MeasVURnkUY26Vx7T
oG/0PgtSe2z5/n2qEUrPHmjnXhKsDh1wIYDLq2zYxtGs51gY99I8l0tVABDbcp8OzA4gV+5r55+U
i+26TfqsS9KjhJ7KqLiuCSnwUxtihxDi2PV8mbpgNdFA8pAwmoez586XVtqYek0601RN7zBaQVgU
r+8Zkc3/3hqmjkN8+yH+NS2RO77jv50Yk76Wt23vmo/EWQj2uBL5ymd3ZjB14e1w9snE1o/lF7KR
rrmnui/SqCk5v2nZVpmfHNi4U9mI7nQW2N/ZHjb0AWHInQjGXSG3ixqzsEpyAZSUzGCveAfwctqw
QyKGwjQzj8OsNvYEfP0Z8CuXxgnwk5f/7lWJdlgehYVgbL4JW5GATFfujVqlCBk2jM7bdYRbpGbe
EhC+Q5726uug0dOniqGeKkNSIMM6pP1X84iOC2NemVIN8DH/UA5o7Tlqg8PTh2AmZplhHNOP0g8t
p6mWMSOa4SQbYgLQXmn9yYCzU7O7HtL1Sdw9Td05+heol4srPkSDU8NGOvTwAFN+M4ax/xYqdnl5
p3tLFasASuURVvVq3tZMcPodcOf4iqd8Rqvb7gdv4681+x0Lr0EmXzMwUjqM0pNJOpmUq0QIDjcX
v76IM+ePZVlB8slu744dfJWfXGr4GvEXpWcmNkG3Nd2Bj/7CFZWuaAsLeliTc5VYUODS+ZLo0BF4
1c9DrFXMyS0XJT0dswWsJx/a9oYXlAX80B9qgX3xL1PJsuO8t26Od1NHG045W7jX4pwtaNLmM9ax
aDw6GVlhf9tQfO5jQEwDIoJxGmSAkE06oa9/vfzwwMztj3f+VP5oHDYLlgB/RmMYTv0O2/lzgfnF
L1xjjNlRqArU+rCo4ANXNBQxrZRqU+55VecGnhbi45Z4YoY8edRlMDNhDV2tkZwYiO5Ond7QuqZs
kLAzrmIX37VNGsppAqu5GLZgOlSv87ewRQtdHR/6Blrh7cZ3bJFKQBjtppq7J4bZuCyOwGVbZ7L1
eQEhLkvwnTMMe1EmzrCTldblTiP1YKYDXAmfPWSsb0XpNVpzNi+P0UKxtQOKu7JW9G0WVuzsWcwt
uumh+uaxriBD9cvxhZGPH0sBu3cRDABfZVK5n5rmFWTAvjIISQmhH0ULoj9ZazmnPsLj8SVl5BPM
2ihesq5IQ6jc9JBxOK1AZq4WvqFlpxbX4wB5aK7ASPcixfqOkSiSixAZS0V5ZeZTSGw/kgSqHA08
2ySMyNPP9i6lwO9fv7rExa9gZjiNFLkF6+x5htupD0gG8/AcEW8a2DZn/yVawkONai5g7zM/pa3I
TaBTvUrUd2DOhjX7dLjxGGRgcXBQWJtwrulUKiRq53Nkz4/9BvsGBQx2EmuqiiQiiCrKC4qUTUnA
uLogJbghMiWOva3Voc87gJnGVH/3+RYD9jIpePQ0IYl9jqEARpMW+sMAnlkbNq0NA/XJj1ptHNH0
iIwonVVd1gc4eJ2pvImt0WDwwMTHppeO+UVU14BFh6pqdgBZg33qvfaIYTMshk071BoCo4g0OUR0
dWdDihpqOQ4SANBo8wNfGTB0SyOW0h2X/E/J0Rts9ONhaKae8C0jM7uVpC/t5QLOFkxWQgNgGl+f
dnKHczW1qtPm+WEeoGTsvA+Oimg9WEZ2B5GTXqExDTp2og8AQFl20K7Y1hgTFKUDNjrZ9LBV/We4
Mnmd3+KEPFtfctXGCjhqFHL8UpeFYSvUMjoPlboiAJc5AuXbZF7Y+X1QlAxyf6nsNGxKdhEnmce8
OSbwnfWNTYIjFwTnR6sbEjKCoWCbEZDO/q1+78nonuGkiP4GdO33U1IHyZiKnAEk+dgb1NNrk3WT
1K+ImGcBVH7IOSodh7Kln2VM5FOubxOwiUFPAowCb+H9oZgc9Cr/Koi0r53L+IiwpkLrLwENGV1/
P7YXc2ZBHPelnlX1eLPEkjlKfCYsPPLFOdPtPiThhZhrW4OmfVyUNx1HB9vVaRAR9geYF0ZTqMJT
60kZbIA6jyI/3ZojRmXNfNrw+Di4Hvrus4xVTNkiBWmbB50Yp2zU9VKsNn8cPolZOz2UWenHBDnE
WDQWXGSuJ5U02GnQrmtEC1DCc9gC5on+fv6Qyn32mW/pCWCRAJvXoZI1dfEyoMZCAMgEvrpL4ane
MD9uobJIDnVPLObjYxqyzoOIRCcBCrpRQshZyYCjdG762oaP2fgVdVKVApz00FdLeYZce5iEcIS7
5eYBosW/Cb/hE6pAV1N4gMAK8fUwvezJTEfvxkt9/xW32qAsQkkPKGAY8Cq+/XpC4Ts33Saom6oW
keIq9INvfTvPPRduDpi0562ut88pQrpiubildyCKYxtx9M821MLBxFJ09G/XUVYoZy4qY4jKUkeq
T4RzOahRMXSfYylDNh3p5OSEe6+WPfLNyER8DswPMR1JG6JOl70Fr90dFiof4EmmISafIVx3xBLs
5MI9WXt4bM9mreHlWV+JycRcaHCVg0oKCqcc+WkbczeUhZi1VTEeKkLp/9ySCIO0OazwhfTkdabB
N8/bi50AY9OXtbEb4IkmIx/gm7VIa4Qxtte/MgNuDBujBXE1K4Zg/bJEHA4Zbcn6k0eSA8tVBkLA
sRV9RX+kSCHySrX/5GR0tta/5u9Pj9f88CtmH9Qr6RfNze78fQaAKkwc92JwJSBmozHLOYoNpXTA
vZqYjjh5eGZkNqjOevIsij+KBaZHYLEw3AdAz0G3vA//aFFujrkV0BHbUhLcLJR53KHM6vmd40GW
kIG4YvM7fz68JDk83EpDSVEk4DQWqdrT6CWLhpPl5aKBex0GdZ1gQPaI2psp6eBfF1zeL0TQKuuI
dlCXeIUjFrtqhs2+TtFZytooJqMfDpK5NKWNxFGu7hUhf0yRk6W20l9BwPnpfhzVLdkzcV8OEQV3
FIAsPYPDZUqjCBMcW8YTFjo8MrD4vHnzSb6L8+aL/OYT4CP+g2kzMoejlaXUnlgel/9VIhDVKdwf
V/xSUwU02AeWJ5RRs39b80ZyV3XrzPtqpwEtfoPxr4Q56jHDCntzqepO0gcsgtRPge1QV1XEXBJv
deMoXG/67C/BSvO2znkkZP3DXAd2v+DeEa78ZdReR73XrB1JLkq21zXmEyOdFrNaJ+PfKCWmAlKk
xFx0qAogNbHDCNrc7c+lK/mxESRcPdTvO/fp8Nb9E5SeN2v0fr/h6fhheNveADdaZbOpiXAwFzhb
rEk1ZIBVrofwz0UIbZuGnQ7yNUzpNzvxoKvqLa6cy4iNFakJdfo0yxVlvg90gx4bGJMxtWmyxLk7
VYa7UKtzIKW+WW/0cDXQtD4g3RHOImnzCALJ4WDhaPRFKQtA4Mcxu21tH1sBOWIXjfe25leWzLhr
CPzs/A6zFWERR4LntEL7kp0AfSsmNZ8yknVdtP5bdp12L6fSv55YPls2dDS9h43xn2Pjf6C02AU+
I3FkQimNdLAbt/pP99El/kK63mXN5FA3FJnaxAwjRnmIMGO3JWjUQjlLAiRKZRJlyy6tPgF6a3XC
MvU1vE/v+luVeEL8qJdTb/itYb4/S2yeuuRxaOvlxGtBA7QoMSjDm4h2xO7x2hkJVX6FaucgZ7x2
G7LNB8pQqa75y3ZvtLajlbX6UcQzFinKLwW/gBAA2dBKp+yhv1ia/UVu3qHXNrKbrYfGuZpmpewF
7aaJxbPVGNqWAcDO545nwrpbNB3Yf+jA4Gmasz/JzPj6ZGEk8TOHVTR3mYU0l67pRjnRunK4FMeG
kW0H43NJHWTRluOQlyGtw+xrU9dFlrHp0Qli6WRkMb36lZdYMmkSD4EzqLf//R0qX1X/Tr2rwjjR
6aPhAtnwCEs/mVjYwkgHQ5mUkB8TNEyMtyT+sg5Wvbd9Gqviy3o7Ux3qDkUag2KInGv4skymzDiO
flQeD40xOYjebocFEanrLpY0X4CltvgdMAy2mmE3/ZxHFX90XXHRED7pIfPyr5394BLKd2Vy+xPZ
7xthf1OqG5cvJM4ouBSi4J54lbIPdFw/QHyKLLl0VlSPwe6tSqYZNIg5SxVwgiiqIvHzVsDzLxul
74xpug8YeIvPmjlGJzoJT9USsRNivQOi10NghULs+K6m0t+FLVthKz1SNFjLkwbDB1q2lnhrRasn
PjaU18xwf50buN4heuPNc0MnDgyS1T9PfTgMPCw5G9OeXoWiPzIEMl31JGUoj7ksG8raXpdH1t0b
BK/Ir14kFjj+Qib3+idOmvwGhO/G+SwpoSNtBkVvFV2yHsufSjhffLshnoLi2eMhoDuItD4ZRoFu
YM1kX8LSSKpCgUEf1BDASLqpjGfiTvhH15y5iA+6u3XlBL57kUIGud3i5xR7xls/EibDd51cZUbe
1M7sCIYGZ/UJA28hqjgpcF+qAPif5UHEXuaxvnOWON5hNika51IYFXZsjWffQpAnnlY6NkKIKfHh
9Sv/Kz9Lpv8MALpPA5X8Qtr420sEiZmjnJMesDYYs07wsDABwvc0UPOBSc7V3TJfbvzJ3GUpzOEe
K2213OblEzscOxfQ6r9beoy/XHO2bU8TX9mQJIxPl9Hdp9seDDv73XBzCsCLq7CppoGlhuge0wYp
1NSSTFbpNO2wnF/NzbZbqGo9beaDpsvBPWii1xWtrJIjTjd6m0mVJsUeQtCefxCC3LIjfggKn41P
dfzKbMR1YZIxS121UAf2FH8JXAftpgMG81v3NEFcUup0Sio1znjYn+FPhnqvyjeYub99FMR7Fzxs
KbkTymA4PejMoCCmnrjuv0u6AzsWrNcLDQqiEcTy34/HCGJOJtD+iegziXt91QQW5RVKu0ryjQ4J
JNudYqvz7wLjNh5yEkcBCSwbpqYGDeZBUYpcCqo3ln4Cnk4VG5kYM+XQ+nm/kgvmf0AZVSywN1B3
N8AyNgN1qpF7RufS/2f9d8p8IcMVBqTTnbVDZlbUnT/Q02r9HqSdOJVoJ04jU/7z6Z9vuVo/tpsV
YpNgyXp3DVTSvTR76w7tFCRbpvQyleygWdXf3jcFbpiT6kXjsCl3VGzsNQW8XtVm07mCOdezFfXb
XmgXXDVdTp3VYZo0/TdAVOru12hxIr/0p2GHI2A4A3ll4dFXDMEud3nWYauXCiLgDqWAUAIqa8WQ
OvYfhp3inpddDTdd4++AouB2tetHR/SOGNahtbKhOnyzdgX+6OTQjPVto+7VFx2U0xlnFHuXIoqD
CeHWn5pDrx1Z8cuqLb73+L81QyyiD/n2fEWnks9xuKbpXqb0fbbZrIP+j3YJWg6IqVvmKtwIqClk
7cqMBPYLX3t0W9rC3347lcirGdRHeNGuVwX2H/PU0CzGR1z85jzfqCRMHTvhWHOZYn6UnR8o2cUV
/64N2WBoNXZAjxSmA6cbq37Vv5QlTYxpwLL+p8lyVCbmc6LBswtPMPE45ggKV7uxQqLKzEW7OGza
k7dkV5qVGoD/JHGheQln2XClIKb51bkcHPhEJqB41a4mHDZng2ENOejnpV4EHc8DLjtfgbrvrCaT
q+B8XH9u6krqys6Rux7WpdO0hSuGxleBf7N9FU3LXqZ6ajoRNYf1zhWupqHrohJfBXE7JqxbLlD/
itUdqNG7cyHtFqk8WdZscxVgZu2ECdxBUekUG6DyxOrZfQ/MrxTQMNhrdHfb5+luQiEo4iNUvrjX
MYCeBW/Ejg0UnQ2N9ycRuCB6LOoOzABHhE0eeRR1TYNSLTYwH0j0V0eFf4MpJzt/eXXXEY3VQzV5
U/cKy7bcbmTAxY08xsfAmRAXwcv1RZCch5aa43umRUPT3QEbph3TdUQkUgbsFKrPSxt9t65QeoV2
u4eQuLsbs46ooMUNhpOwQwiDnirVUrs/LEoKGkcg67TO9qrv23xquAomYXbfO83Yr6qpWzuRKt5+
JxViqM0GRCvIbzxr1DJMJP2qqTURpbEq4q6W1HMHPPU6T74gUgWqGC2Cd8OBTJ7fRc1Bgth2TMWy
oMldSgwD+AuXTKT7n7r66He3ruwHi52PVKN+sDhF+ZdTtmyXb2OkOEovtb04WTbasrFcybp0+nr/
pvlOXNmVgLnHSkUUd/ydvvw69taGlRJ2SFR4/M7oy9hoit6PPVVb+W4+DvbTt9++jEfFtq95ddwy
RctyZeVimScu6wa4ibzsXAcdqUccF0nXSspS67mAKIlGBLHO9qKguWp5JbqymJCIkHVpQcIMu29w
jfV3GECK8//O4+HhRqd93iKxGySe4jAhXPEk5norsA5UlBAKXy6FumjNwuo6c/4mSCGMiVZ/4icJ
VAbqVI1cdUOVuhW9x9e5s98GqbNW1Qd6RCwKU5cXZVPb6nWeBbCkJovDKmyOtHXxwoTeLazXUiZe
iTlms89O/hypnkyB4dFiwsOqgUD15Smwls46r3aDVi+dKNGCIz305YQH945KWXlXfcLMsbYnGdtO
8L3NYUktOBUNVFKZjvAT8rB2hBfozPTf1oU8+zZ37sVBG7IybZ4JIukYdJNOYuBCV703uiSc+WI6
+ueDLNrIjSle52RCYNz5Fj+S2MKdb5M67ZmP1JvsZrUezTZGa9LOItNN7HhrhybCkQ1wC5+ZVm2O
A85bmOi9qkze7ujt5g+VxyPFd275KghoeFsCTX3UVrk9oiWvFjM1UHDb+zjjVMJohFopJUDxQbUH
dB3f5twXM3UCTeEYh6FtkcduQXAm0sSolO9nCx1/PDSM1O4ety71HY1b0lsbhx0X8tkdvBiEHI3d
PM0/9vIdrLJzO7IVsQk5bO8GenAcmmhGBzeXaYss7ymJ907k7IXpXcVO41dbZiuM1Et++gOQR1ZA
WYdiFAUFy6o5JGm0TXg35YfMGrTQW42ng5Bl2jUMnkK5T8u8hkeCQEo8JQtd3l2rlQHS+wLYktg0
S+rorz4lSdnOHcwdh4WYQOQDAEkUinaCWDkSYcrMqQAvMN+fORNrHgpa3XSkWfAVneXnY2OCd51y
B05tsIT4Hpedum427LpR6gB6VS5CobUUu+8IhE5b3AV92n3ln00qp6UApCnmQR5jUCd7SAewXmiE
eaDWhjvd1CvBd2rkq7X1dUygwkRnSmv2iPn11CVTS0nRQM/ZcX9xxmnF+XyWSyWHhNHB7tURAaDx
ct+D/7nN1C9Mq+tRIwksaZrO4u8oc2wfLqp+3H3NNG8lKSHE1KseMMtUZgMlTruya0+6cybdOETd
GOJw3P6f/776OonMfY8KipX8qlw3IBUtn7O7swPRwNwb6aOx95O6EmQdVxN8nZU+OigpK7A9EaHY
pMTQPZuJpZ211REmmHL4lUwmbt5vDPU4x1kuv0UlTK9vnm05KvcATTEPvtb2a7dfk58d3jYqHCuX
PIu/PkDGeECmC6p/yDrm+qBjh+X7oswa7vL+O+xkh2B9QMyfEkTYDCCBa1qnW67d+uYJ3pbKdMyh
74Bc4xVtVfQuzMzoEqIvH3MYCvOeVaNNMA3vDRX2dMYI9Nf9+cObOnEvGRMETUelbwNWXoeGkD7E
3oMCy0OYu5wXEbP0xDUSBKPiyjiPpT9GFDUfhbuHUNY03eOhvaJgnWkIC0rE+5qUBAs48+2FOltN
O19yaEBTCJj7gFZvPE8T9+H6kdnzI9yimHNfmYER05ZqH5tN8EUEEN0BkEp8qu4Rf0M8IkKxyiHv
jTm2csXsbrklk10XZK08vN9SUEBlBbTkIOux3QdRES6LvGF2ykJOg6glXGPnopXn+9ecu4boBNph
rTHhHGLeYH+l2w8xRbtFta91gxyPQXgV4+e5W/8JuMaXcoBbgrLp0AHCZwnVM9NaK12/UAUowhBG
qC4mBzHXWQ4fE+HuMIcFgcsimc8XKyIWDmrmucjHUJAtDCNK1lLh2VyEfZlz6YWRFVOLpoygXxyP
iNTI5358DFem8WxPNnMOyNb1g1dB/fmwkcp7QMJFAOJBjJhW8KIpn0qHkQTHR+AaqF9vJ6D5uYlJ
QFruh8LgDdTcW15Dh9qKtECvVlsDATF5BAb0lQAndtJ2ULF7cNeyHtkuRqxG3yXh8agd33o/qY/A
7fIP6lM3XlsYEfrBlGABKsKIhQDyuUE5xLJYC/inMAeTKA521+r9DBo2+UDYq0JThozSghQATs0G
ghcm/NJD1S1evFaNGWbtALz9vThnvITSaxSyaxraerWT7/XHN3YG8NcTYitPZWXREBLogn/r8Qck
lAK/Re9XgbmscmcD1+486fwLQNu0aZKanmm7ojC8qTxeZSL1lXm78aVwgUbEhfz7ZfOa0oBzstC5
ZhpXZJ+iEzrWznwk4GM5vyt8DnyACBChqWpZR7Qwr1tEL0YHjVQ0lz6PpOlk6yGe1CNZcEBt8R+W
YUKhkstxY5/1ybSOJJBt01WRgQevSHKUuBEeKzupXCwS/P0DYfzkkgieYywZEEMq6emBn+rLoBx3
NZy47JqWllDHm3ldxiA4QNopwBs77/Y3BOZGlZan3UIFkYPG2ruBn2QZKkUC7lwRAwF4UMFL03cq
AW28fJz1FsO88epuupXLrkTsMn5CzeyvJQh7l2hnlm9wTLBeQ3JRKa210KbA/ImV9tJIXaV5EAVl
EYnVXV6V3jWMHso5t2SKM7tQ9ox7NhmF8IbSFVdje/ZdeGTSWXCqBi79H5Mqt5AOBs4myeYo/8NG
MUgjdcCf3R6jv2mmCf8T/xP69Gc+8jlgKsAJF3usj+zvFeLIcRIyUZDP5ZMWvYYFjBSkoq0vJcZP
46F6l+o3U1FWA8FQ02zye7b69GF+DjRkW95gQv0CHf320YjulP64GRhY798h+/iEZFUuHykF557d
NBvfBzSrJFj3q/6wua+Nzv0nBfY061LsumSh5E9yGfIWNakaV8M06wVchoBY4V9hkWPhjlUN/uBq
s5md4EkoyqA6dp6sp5O1rWOzq9OiTNBqlnzWp8Y4jMk+rY2yaK6K8elbis6XUoXdHa6rtQP5Dreu
W8i0Qgysc/SuAh434ETHNmpS92aT7tPXuOHw7kyK0c4fHgxhvqyzVY++OdSuapU6wAMTcnE8OJe4
QBpHuj0CauHVQ6QPkcFXeD2UQRXctoaR4N0+6gFHoY3+Wc2yGiiQrBvtPpsBUVM73lwTulmfUMUl
V2po1Aqb4ezz1xFm+Zz7ZIIH0PGgVcSGKW6f3XEClUwzUVfdDstFremIg+Mdp5xnchLUs2ugsvIX
psZgru0omrM1oTdbxij6OZ+/fenZzdC0BvqBXl1Kh0tGoxMff3UgFUiy4dEOOeCW4FzMAYSaK4EI
R4n4Hd54kF6aRNjeWIMxzQbUMLaPW8ygpQs6y19S2CbejaPpwlhkicjhhhbbRO4/JQzdaTb9goGG
J2mcaw0/DjDBJx4awwvLP5CwtjWy2bT5W4hrMwaF7R252nSYc4yVlVfTsQ1HcDeQf0FTmTIibofx
SHf6OvudGktfxJxTOSD9n92ZdLKMtOZebUgENRo3NJS8yaV9HJJyukx/q77eHppYDv51qnUgSHsQ
pRtshCB1f9XPxz+ULm/HsvpR1YMc45XChZPTiemnJjxwKjZHbss0b9VXk0Kh5UBftPPnLXUn7PbC
R3CTdKt+Ssv4H/DkhmpMRvFPLyZ7Tt7e4pS9r0M2yLY1DKNzm3eW2R/5QUM11tzxtnXu6m8KxdN5
qnF0Xa/EsOn/c6MrrVxIirdVNMNsVWDY26zp4NHTGE6fCN6SKGl4kyApNcoOHWCu0vVaY5XSF4DP
acMQrOnN8N6WuVTtG0FCgHgtqsCtlwrtGMyyRUe9SbY3lim1CRCaGK3iLNo/DvyNIpWIJqCciLZk
jqjUy3u9iTtATYOL6rnAOq4GwhlZMMhSzU0DNlsNzXO5NIUujceKh4nqyFBmBGsyxXIZTveK9JUc
3z4jZsqdobpP61tmifi0VcgW0mNQHnaa1rDPglbFKP0A/0FGuyT8N0BogzbOAvaevg+F6jlEHdTV
ZwlHS1vXSHR55iF7qrI6AHLPW4R2/7+EF/5a/4m5dRZaUfJBGlInoiAVL5uAGj3ksEXYUBAko+yV
PvbdJyqVMkPN0XdWoVTpTRs4fCDHqyyVSHXZOuGm+KLv5x4wc7FVANUUU9kXYoaGZwi/uU+9M+Hs
C8z6TBrBqKumfBY5a6tumv3hLEySeI1Am2YxXdSkNXCLzltYllgP8kIzRrBIPUegJirN2gbhngEZ
FjJm9aeyp8kVP9G3VYawPQnrl9Ye8z73BiGklXox5gyWan7q/Y7RQS22bEk4rfZknEI4s7zXsUt7
GZzTjeMxvvRXriEEWWTbQT5zbRVdblhSzHBJPhPWqhTxqcHMCcsfuxCH+brrwGsUcn/HIhJWnGmt
AJ9aXQyvaZ282FDQyUU9sQKRLI78SXQcLHx359aYiA3+8+k6qYcjOQdOTnyFF/VRlr4+i2uVQhP2
TzLulzL8+S2I7PcFPCeLliZzSBDC4upO+AztGJ1XGrxhe3QvSQodg70UnuSxtUcyvGn7hnnfciXN
m+AsiVb4s5jp3kxoEuzkvGIyZ8KGklhxpdw+tvjtWKBBg8B71pQa1ZQ5M9A08q4MWKMk2uR/VzYj
JkNutSEmuJo9Lbi7f0F75d+40bUcG3pxfRpKSEe8SWA/hh01zU1FzHj8cdYnBRbhV7pLAum8KoHS
TkRXkE7K1tPzZdN9hMYyFiokMFw+uwSV6zpYLn+kSl/xP6HACGFERxzGNZWkIUT3SXgAfVNsRAvU
Bm8sB70labB+K1QWXlpo93tOgQxtnebuM6Fd+NUqDw7lZa8HkYRHct+QareME5kRFKMkvKO15GHZ
sutU3kZxwl4dV4lZD5rgvEYdxzwwsMQKeFl6YMxO7PUITMtCyFTzZWXsB1wQ1rGs7jQfCr5aqrh8
VEiOxIRGzd352iZsN7Jfao+4j8b+yZEmKiQq3rRdLjoiRyQy8iq1KxK652FEXBYoUTp1tG6nFyd4
wyXb3ZoqzKNmKSRtBLOt4/rdYuSpEdtpSPJK7CeGhI5TVOxSn/AcCALk5HVo53JLQ9cNfc2IihU8
wKcZK6rT7xDInw03T87QdY7gX/ofxwOjyzeuGGxrnaQdQphUL7+c+c0BieYB4beFeC0GUZrklRoT
zgeHt2wrWaquuksJBLJHfpwXdF+4+88sVsPz2H8itktcsh84AO0FUb8D1g/pfVnP8Q0ahdWbKQ5d
fHQy2KcXSlBys9BH8dU2swv4ZZ6bTt9cQLfDdKIkR5zZ50ZqUpJ+KZWoPKDVcsbThusRyzeFB0+Y
qQL36ZUTuJqNsC5xD2k9PQAE7Ixcr3PXP3khgeqNOWwAAxRlxv2uuu9Q3Zmuw1xH1hXMrPP1kLXq
n5saHwMf6/UEuHEoMGrC1/TVZvDJqvdPiWPsiT5vipDzM6nOQwo/NVx/jXRvlE8ZO1LO/w1hmRoS
o8ZGdv1CPuukPNqRixh/815IuXv9fiUcz5hg334A24EK+VONIokbVlwVNyrxGgHUKdvJYW4DR+jq
7udJvsNPSY+FmiyiIH9ROFDDHVVE3nS5hDIk+CwoRp7xo0wb9KTr/KcK1so09ds5Zdt+0Bm7UOQA
YgY8wO3gyysGe/XhcWRlPS2Aach01aFOxzL5BLUJkUqVOQCIsZZv4UKIWaiJopjTsk0Qg8EYRqYI
ImVQm+9l8rcspnYGNtSOUe6llkWn4xr2pfIFUZ4tl26i5Gv61fGsomrOOHZRSsaVc8vzKKY8siHK
LK7QP3eaRgjboaFazJy25CGi7hqWjWVXMJyjfse9Cea/5R4UctZ/PtOMag2ej5fVyMhnCW5/m8bx
cQF3e4Hqsuy9pqGPcJb6quoIrKOamXOVP/8yJvaOm/P7Hj1IhCup2AG49ljHMEa1MXA99v22Hsey
v8h6Q8qgIJwokcK4o+Kw+Si10UMSgkOoSa83e7y69mA9f0kR+qH6LXMY/JkkccFB99gws+9TLeXN
GoV3b3LKfK9xBhV9PWk4h312JPvI0XqacYoUZW9O2OO2LtrHy+3GMZCpAQzDTOSQnnnxV0YM4oPo
yRbBk97MAtq/69tW9bOdqAxRXA20agdEe52ocX6thoBGZOjIMIbFD7h0re81fzgsJvxDDxDnZgRT
y9qQI42AZXQLFUZ532T1x5+i6M/AWTZfLLdmP3oYKE1vbsDgBQCbDvoQPSMcEj/XXBmAWizhW31r
4INC6pWvbw9v6jNBy2Qzf3HMnYZ/gi3MDyUJ8oqdtC9pPswVBb61BR/f0blzPDJM9LEHejRyepxG
W2OX5dYXqQhDyJq5EeBnMbVP9pRzFsvqwJM3gHOHxT5OgtEco4RC6c4Pv9s+Nq7gwKB9m7EoZP1z
NtxO3KOk5kn6ZnJNVoBb4y2OCSopMbTWCmiKMh1FBSrpbvirla16FNbWfbYHiDvqprUR4Hqf39ES
wF1fIolYwFMz8p39pz2ExymYOPvnDa2md6e2pP2t4EiZHgn987mq524dePhOsbRHFJy/6B+kSJ0F
pf139DzlXUxxedD9jMfNRgLUI5IAw1BP5MNrpzVHFftx2UJVrEUpVO9uwXXP4hFQT95mAeS6JFCn
bj8Hmr6cWhu1ZbaDOZLl7NRPJhvVDESd35NTeIbk2xhxEhX0mcm9LwWGCKY9NcGLojaa0aaYuuB4
Msm8eMx1QkgYAAwiraTQE9CbF88IBC3eK+ZxrZ8oPmvl67WFsJkK7B5/W1b0S9Mj3fX5WVWo7KeG
oHVagltlXZTfl86nPZXhDJogazuxxPbcrmeKkQf5vZl9A04RkfwxOZRPKY/FMutlZjU13Zl4yMA7
7g0K4AsK8XtIkjjGj4ZZwakfJKGsojFZ2aydUdSvEUAT2gzTETuzdX0LTVvyEEPPaPz2CGOCKtFb
UzDKQ42dDcklnsDof+dL+GDkSavXhDxUJZxVYPvGDu4PBqb7kMJqQd+22NDmBibNQ+0w7EXvra25
nZ3a3bbW63c2jA8p+G3+kPAdKKLcpU6/91N+qibQXAUDva7g2/8TvXuuw7qe7j+ylJjbs1q/rNnl
wk8GhgfFoglknCtvXSWacf9tHR32525WwLfC8QAJ9+boPrT0AmV4h/g+wKtzJfu2s0QYjrrg39bq
Zb5u5ny5IUo4bqav1DnPcJq7Etazr3if5TPdzBM8uiykKimqmnJ5Uq3AOf3X9QiM8wRYur+6KDTr
MJlo97JYkpPmwWM1CSFfqtp9yJgaFVTxiJKjXLbm/7AmKYzSKmfIeTiRXQpb+hpzV9RnDyV4b58U
SQFBTV0YkgGoj36f8PZRtQQhQbMlsQWIJeNzF4U5sHIbvM5SkeYj2RM93wVBypugVvyZf9NpoH+M
XTk4wiIKG9KFooA4G4eD8MiruiEPcoaRRdOwV7OuC6OZkPVatjxAbD8eSaxaZHWvql8wMXh5o6T/
kedDQB9cw4demwpcSnwmjmONlaAmSBgWcS0XWz7FgpOWjybz+gqw4mv3T3dx5jSalIv9LJWFJGm5
ZsNMknTFnDiaXvoqvtSz/g1ccQnn+qJmxau/MdKOGbELzHLoBUsqu18BSGgeVZn4GqAK2V6lGcNx
MHaHLD3d0A5SAzFBMdBhfAqyNNHvev5OnG0qVuVVlTs1MrQWAzmIFujvbEysqwTRiME2egNMZYvs
v3QYxTvYbwo2YkE0c/GXevq5wBt5ukn5fZUCEJKvHDdUHQiaSSV7wOFW+BGYCalCf8z2EcuCaMy8
7z1nTxjyePhZETeFIajfwqFZx0Guc/1zCIf7twXl30/oXKSvnO0KRUpZ2TWdgjZA/R7ZvK9o6E22
L1iTiMVK0IQfekQS99X2o8tAHen4HEefnS0x21rwpxIKJ3CIfekIX0LQ4tPuUUCM9nPg9LGqZLBT
olWqZliY7gWV3Xk5OkhuoBpDJZYpc5Ah2iHR9PU2LQxzk6kPkpeC2axV17HeAWfxaBTwx6on837F
luqLwFbQq2KMAqVO3635zkhegK5HlcxCyGTRHX+Gj4fLOClk34NEGEmqQnhsdkMGfa6RAGoaarXK
UHvXR3T8rbXEyZtQni4fhE0XCri8QuE6FsHHPJmJhP3FQnmlcyFITpxx2fxD2GuYHq7PlsVCyV2X
kZQ3mQ/49xl14KbJ1gcBsazm091dIHW1j66I19gf8/JgaH+9ZUEVEypbUvrtzPShOCKGlsC1R6PX
gv+icd1N7URjkIdhsYaOJbbO86VNg5GbWLruz3BDz5s7SYBtxGgNY1wCiNscb14Exe4xUw2/ZD0Y
ZgUFE/4/E4nTHsAGWcT5gP1zoB5kgubYUa2MALue24Yb7H5vCMkpr6tWDaKJW3jDPR1uVl0yKjXh
EK+SK6JgYhrwVj2fN9gDZkyU7FReFz12px2D9rhfwS3VquzVRr67fzMC2WFt0W/hOZCUAfLEwss2
YPcojGkvMX+iasX5ZCy7eLbi8nPzwquugXxk2eKbCldK0VgubZNfzWopuCEiQ+VZJHenqAf+hhpJ
ruTY0c0zLlFyCYYxBIyzqR508v9lHbYeUKKcnwKWAmYZqdbk7/KoTeXvPLbPUkqCH7ZNTyCguYNA
Fxjr/72GIpuT4PLHLzjFVlaMgaVTOB2o4BZwnYRdASVr/h5T/OlXPCrdL5Tzpp4gSTf1P1gw+GsV
NBDDyZW1kY9rMUqTEdYuB91slNOPZUXBumPAnPaAQ9EOL1BC3mEfM9zcPaNSZIRpSq9SFP6q2A7i
UXqnms+8lmK1s/lXF+stibT9SdVI8al+7D4OfQ6+qDuN9JMyT3+OJnZCTf53ewOrVRSbMyGwhCQa
6pFo1rKSzoESsiMVnN+GrltJSKe+Btasulal8PVIHBS5S2kwWUCbsUQYSq6BDtv5eBfJkIsvEoKy
2fTWqvzP1+JJ9nyNLyQIDJQQeODmU8f4NCQEKeZ+WW5bqZrXRLnPA1ILQdclVO5M52o+WD+2qvTv
+agBlIAlcbO6Tfv3h8OwaXc5cr+DqwA5ByTjpsn1Ie1IreBkFeBLZ2Ak9cWu7DhoWVqZPGROwtpg
Q/iWN/qf6M7WSKVDuLDN650+UpYkSTm3X35jfKyqn+rIDHDFjoqzMW+Mexa5dkZ3sm0qiblY6cBI
w+wbpj3yO2BR6WcmkcYD9ZUjQm59jwn3/wX4QboWxKKw3bwoLEcFjweQelOG3svtxvUHhUN5lnsT
utmnNsViH8j6BwTOHuPU/s+E/XK0KmjWdUMGDYg1fmbPkQM9P360raLvP4k3WY6gncy+8lBtC/4f
OjhwOIkX3REnuAYxALBLkYaaH+QLxGFtewHL3jEjXtBeHwOwHCfZNnn2WnKgU4Qye5RF/ziCKVp6
/dNqJaY8Riz2KuYWx0SD6LXTnhqHmL76zVpqYadtIDlg4BUl8HgXZx4OFt7GiQv+s43WaAuVkVZe
9ZXKmfXBenddov2/T82diM9M9itWgff0rhUz+j5UGxFuwOq0d3XYZxv5EQvAMzFc0SWox1/Wo02P
9zR2jOSZpzwvdHU+3ZXbRscS5XYOCIsKxRryP+BpfzioZTbDVdXmMvAnqj3ZW+5J91rEEi47SAVX
1NeRzvY1NhuZAZQTQo7gM+Bg2uB4Knv/CpfyghTPxuHgGNxkoxaR8vLboQ4/Zb1SOVzuxnHoaZAp
5C7Zkdkw/Bv/ly2LUDcoGiG5lWAtRWLzIB+9MmDl/3ByQyJtfROVuMjATF0VzDHfclOPuI40I620
rhtiV0winNxg39T8VFLosaO2u3duWmXQD95RuLYiFh7quJbPDNkweGFm66YCo6Q9JZnUkm30vJpH
OGqPLX0EUhOb2dSiDc2mJ1ZGF+y0EMswnHuAxnNBqbVLzS3oMPJX27brpwfDtD6tDsuMIGKGssBv
K91niMvIkiUapPhO4GOPj3rQyyBOlAd34kTX0a+3sAK5ix9yjUONlG21Ys7H7Oc/r49K0coHCWis
abxJmLiH4AJihaE9h1xjlCQJNeTUKAzRpgnQ0FNV7+P45bQNePSFJpGMq3Auzc1Ec/o+nNpIQFU4
qxmpMVzZQlsGGTXyKlo9/eDqExd+3UjBZZ6siqPyOWkukvikqvkcwaIMX6DOBYr6KswQJIC4WNWw
fTJT1Tsjrt3sfo2Mrl9XvJXbjV+AkaU6Sroh4fVFPtwzM4QHL2YeqOKwb5v4Z6ylZJ4n9Y+0ywFA
UO4cqnIgkFAfzQW5R+kgMlsq33Mjf3k0z+VWk/cxW6ubDbP/vVPAtLszJLdx4Jk1GqtmbPWWU/Lz
88D8X+5d40M4mJljIvF2GNrKPhKnJMLEa04IjV032JOKh4tyrgLhljoqtXBTC00tdUD69OQUv99Z
U1+LODMuJKZkTkzh1pl0i5pfWEyCzqCYW+95l9MLq07tz56sWdmXPxUSrYgbf6Xr/p6n9pycbtoT
ZGddFPEhiGqKTOt1Za+V+6Yx7gLXVwiKr20sOmml7KA2mY+51xLZB/erAgRPUKYDEPEdUQW01Hvk
k2BNXWpb6uNeTmap+AfWxoSi6suWjT+QTmrFwHhbSbj591H2e5OGRYkcsCoUsC61gwBlWObQH2iC
AMBhME6TV2wOCsIdP6gKbZsuXN7KGAJXXU1PS1Sn6QzvddzFChRhkykID8jxtYOl4kzZQWk2XJhy
zFo6pDbQ4kDWw0MUfoLL4HlW5snZwb+ouUXpYkPCya/me+rX2U2Mn05iF6B1ERTpT+R/d5fJl86z
0JhSpZEzM1kQoe5hU5Xo5+Sgl045d6MFjP8MQU3dbo3ii6XEwNuJM2AOMZeAssqG2OxVK9YEq7AV
MW3JoSIw8EIDHsHhRNYY60C8DV1uYp7h728sOsjLuHfgyKlVHovMtZGdfcblHuu8VPdl+1srPdtn
YPQVPc2vPuDQDk6Gd/vIzCe1uFpIrW6NVgwfIXwncnRU+mgH9DoP6oic3ARGVMiy7viV4YqJBRyJ
fN8a5CI5XZkbV/3TT8vstAfFZSsY/q9THRleaMjnyVMAOr1N70AFRzLbEEbvc1aRh6ImYrg9Pyd/
PCUF3hiBODvCeX61PxAoiT87HXAoLI6xDVg4AZwUObiPL8J66Aym7PTdn4tp5a238YQ+G+iF/4mB
TckmlAeZOM/F4q/WHOTXGGUkFdfe0luLEW/KGgSHLMNfQsAwjyxdniqjTAPkxY1hTZy0mzrHwI4A
uGAWzohNcFnvxnCW7Lq88qbIcOThwWs6vXtHm3iHDKdmF2w97govwe/rcobbt95w5Q5fWfsUJMh0
3fkKpglL8/sGai0uOmW7tF02pvb1PZ6cYOmkRmJFfGggOmyIHmeWjNSY3ZKpgS1y80AfZJL2R35d
5NVs08Gs5xvDoTYdwKKnXus9LFMT2Vn3QyUl+w3jgAcsNZgc/3FtQzsvlrFfDV30QdHGHjl3xElU
QhRe6z1/3rnXrHErjlOxgU4j54P6uxLQyH5tLVfSd/vrL4+ULm9x02A4qcHbdzJ7gCrYqynHF/Sa
Zzo1P+PkwOiLFOfDF4CexaYcTVGxIkN/FkihVegMnQd/HSfbDTNCHnnnpwlsPdJAvePgTqDdDqvH
BnIfHWQNUm1921/9r9v7vMZ1a2AIUfm0n/DYUiL18Wyuj3N81Tisb3gdyUmSDG7719Rz7w1gF4kQ
+p8+7kjD10cx9iATw7yE0xphtLEzSOTdAFliV3tztNNFh/mRGCV7lzTP5gphVeNP5wDAhahskeil
NV/1co1mgNcVSHazxbAiXpCS7kI8Kh/nKv+PF+VvlZJJT1g+lOARVRUDlZM7Zk4RxtFr1jELPTel
SnMlSDe/L9YE+SQRMI0jk68LRtGX70MavknpqCGaB+eVYOsXEl103uumbnDc0pEy6QtdVYnaRw+7
UaaKzMpnDVmhU6AcdZl7NldfKMJtd7xA4Zgl52Qval7j7yDtmtPKwAwB+WzG5f/p3o/ulZ/o03TN
PXowKw4xb3hhFLEnRKyqQZNq+WCY7YkG/7Cihs2+iXGm1YuQ50OIieq69roc3211UIkCduIoOK9r
31DtpCxULd20mHiS5Nhufgseh1VWjQeDq4DeCWJNIB5cSOVlzqrOmHLWzxi3XLj732tiJEi4AoFx
xmFAj31jTNAYCl2mBm/Bt8BX21ZnV9SvTU+PAEgpK8vj8xLKBVhQsKzCvAXSqYgeYB85EjrfmBFi
f5vk281koDRdnd6WHSgiqP7p2j9Fpor0V8/I4QFfrs3KVMddcaMzUEvwk0covIjmjuEqusrNVdQy
Uafr1FkVaee6/ASKd4swpDeTdqYDJ6orgT6ZgjqrdLEdl5eTDHi2BLwLVmyHHH/8y6UiOglQ7zRi
7h/R7vuegsjRVZVaHzpffrMaBjB0IKLCRNZ9MbDRmoLITeUlfL+voVwdKVVyT6zsuQ5FPhKpV+or
rHzNnhUgQOAUyZQetOgtiBb5WwgTMMuLGgESlrGxDq+G4d3fy3/dsnVJTAZoWgGFgkustUcaqLLb
Vll2z8OGkmUnudvXymjBhHgouCPbi16Kmk3rH99HEnkXDxoHWTuANzUzx/jJz7NyRum9Z6cp+b7w
xMaflxNCC+gNeFepOlUt51eChPQ1Z1EHYtLyW/SckSvxQZFiaa4H+Vl1SjHKnM3ng1JsJnl/Ef7r
UTBrbTbTGOFohNZkN06LR6gZ1hqS9SVtuKKNUgqRYN2nnp1CbalKpllBlzTbIZ4jyMRRq53IEoVf
XQxktVkyf422AFhpEbf9CGCMS1NskQC8Y7HMwh4yMyF5rtdGKLP+R4BdHS8aaemfQASLBNcCINy/
/eyycKoas67jGGQ6myLIf/r7dzWanwGAX9vF3Cf5h533HFAenudo+mpeA18VFqnbPoRrG3CGYH10
VkY7p3T8VNGEmWCsR97nrLq7AdrPwhg87mWnfRByTTzoWssQukftLtAg+bkPIe4MY2QuzwsUQSEN
KFm4glvdAjxwpz4Nqk2Sjx/vdx6NAZ/RtUQkqrLizVvN+NCwhsgkrhEITziKhvNelOLPmQOp6+hF
8U1RtYuDitxOYqMeqlkNALCZnP22OOwSCEqcX+oLYqzWPQTE0E2WjCFiCCtZ0iQbCjFtXM2qtA4R
2foqgc7zRlFIRbHSV4iCgFCbYH1ubiv1ggKTbHfSY5VKE7yvPDlStyRKgid3L0Wqr9EKDcD3wMPQ
ZqSfLy5L8RY+dJN76SVMlhi9MpBw5Uu5I0btnfBVKUs4ilpGDmHzHTkDmfFXIFSWYkwDSt4/Z2z+
p2EHxdMTr28Seg30CEO9Kfxnl9zALmCw6owg1RBcz3Mw7Dqj4jchic+mmLsRqTkaUv4ndXEfA8u0
zWOOx/EUSMUpEvNjqEvI7lmHsdQqPko96mK7MOFQTOxZJI65KkSaF7oFrZ4DLiWcZl71bFrl21qM
X/uAO3g7jpgAmB9G9FKOnKcIzTE7H79xMDeq20HmAhfww2okcOWBgkzOeudX+bnjIPR/l6Ub5doB
BUlSqfp4MTbEPWvXE4F7urUHKZ4AzrbE/JnyYmwVJDjFoO0Lt83JH0iTRU815z79kCPLSOm5kAhI
UxBCckGLgyI2OHwmLIVC9tkQGRuHvRFSdKaty42UXaowJY6yeetOYOv7GN5AW5Aum9XGpzUVaEm8
dfXEEUx4XeOET+n52eiD+ilzVwjyMhHCCEMBseuC3T7ciDkZxP/SVs0OC/pN3uR3HipCvoCWuw1f
UwluS0Aj5O65KhvV/wcytCfyiRPdNseUp6Ub3EAA+o0qS2wCHnNRyjI1BXpJ1crZtp2qTWMLA4iB
xGW1IeY9d9lSYEmmKkDt5gSRwyMPCVi7V1Q5ANYSvM9+N2TTI2YrqP8+77JN+fcR1p58DLfbaBZj
2ovwDqXZKJKNwMoNSRSn1qaQVe/COla5WP5m7UjTt3l3abjq/tEfulm8iXmkKmB0fjTg9NFbtZjk
0eCTgd+OoNTdkabS4CLNaJuXqEayuUHYz/nTySc7e1SeeFUrLXtqnV8woHoiYnJUmgJ0JTDAq2g1
KYU39lEUzEBZNZGyXdSjpSaeIjYChhOKpe7oku1aexzQaXEm4W833FMvs6ClJxV9tIrjRi6Hosbh
vSs3ty2wy9vcOV2C6iHqS/ZVOPKe64NTIGDZDPmSig6GgIn1T5fYO0INfIgSE/O4k7I54er3Qdby
IPkNdTnl/IkLgPcLrTtUamEPG2TkB38YWwl4Nkyx5uu7brR2MOz1lb3oBvn9NcSrZwzkIS7rPkz+
0PloztDyyp7EMutC9nUxGAFP7o1qzSd1kZqwKjIswjwr9qbvBTFuVTJOjAQ1ol9J8zMTZXzHrTcC
702KNgX9AYdAmw0pazAgTEvQU+/faqRX6/4K8YzeGNLyk2xz0JXU8kM+WlaEcrzoJbOxPLTfG9NW
siMNcso4VNZqfU+WgfPhqi4nSYPtn180hp/+nybeIq6N2ZjrbucSeeeuwfqFoRgDUnYVQ7QVNp0Q
LOQSK9QthmTug3SA8QHpVQukj8s4WEX4Sr8h0HtoWLdE1K1+f+zORJbU/z2PseSoapXMszyabMif
SP5pB+9Gk89pxjjKPB73SJf9ve5cx0tw96NxI7NAuRVca7Jx8ZFEh/D0seTT5M5BZfXYpfJpixRL
wmpAKITQ//AanSHC+jY+tn5SBFQfh9yFKV5DgACWkt/IQ4Ykk75A7MlO/Xxi21HVAUyc8+hzr6ur
bWafcB5VZxHDBFY9j2wWph+p/9ZqWcCCiUJW42IGXM5RoozofJBfN35l53KsuBXYjh1xdqbdO5YQ
cSMy6SBsU3B2+dYYQO33+oQeZZkIRsYwhhMWr8yrJpHOO1GLK8h3tFjTC++ZBUM0o46mHnFVSNQk
gfp7ntvJRrwdCdifEmP8ZilPdQois/pg+MeFY2g/v2Myc7unGWPRIhpEp2215AwQLPEgOoY5WFCE
cVVsa+nAxi+qerFmXrihVVtRovdE07J4IrmkgKCwVx2ZPV3mSI1xXE0lTsYlYa73/VlhGDDOXgSC
oI9T7EeJKBlzvPquKCrBg/9opRNrq3//ys0BkZqfcCaXQniN7tmacsltmcEqJ8T1uBRzrJ9lLl5b
z6inLSULgg0p02En98piYUjmurbpSbcK01XpuvamRqEAkRfAHG71o3hcpRiZiDKOZhRxV+he2+zf
Zgc6Apzqk1VwD8eVwMd4CWvVeVYS8QOmecG3s2iCntbcMy8X4Gx4r5G1Ty2FSu+ZmO7F2Z3ggU0j
BV29ORPu02w/ow5I+rbqc3/4jr/B8vtLpqdcuoVkv+F88G3KwOERGUKNfdYahZK9eTN1qf2GvT+4
srBtqNdrp5gFPDMIK3gksdi4eAg9h7YUQoYLCOQEqt1Lk9EBJ9GNuwVjpTnDdEHP2NMHMHbw6HLG
MhxctaZTrSN5sJJtiiEAgBIJiuiV5Q8ePNOtvDpFE4PNAN7hgIAYK+PHPIJuIQmcRMUzZlODFJIs
Yzvmh0s1mqhvwEq1Hl1RbUYQ031VecswwPTbPzaokUtzQrJYhLtwkgAANeV5yoTYm2T4GuRkxHt1
zahcPaqxWNgcBbLtMqn/QJjy7xhxmLt0ktxfftVw9d9YPgVK2CXlsJTuq4LeH7kJVYPwX9fQl2Py
ogv0JUoEQ4+Xm2YL9X1EeS2E9kZvbor4aKC4iEEAr1joIEkrXnNyVtZ02FrrWocagn+vUirXJw6Y
xFVApeDDYAdgBoLOGUmIfvsf1JbppSMNCSirP5aiH5d4uxYo+z5QqPNIfs3AeBMZG5qhZSPgudI4
eMKcVvBvVEyYI72tC8lOvfYtikGVRBL+qykRxnfJ0D16CDg6WLt/arnRK+5ZKCqPiksHPzYjBNJL
prcVA0iMvl6SxDEb8IeQZCeAZKgtqqM+2Dw33w4mA976pUV72Cu55fR5ONC9q5XQ83oflotjhexo
TULLCTKrva4IwFnPgzMM1P6ojJ/mKf5EdL/jJnVagwAg1pvmg9kJni7jAvaJyGRRsbBFW5LL3Q5Z
XxzqIIP2Bk5pegb1v89sz5Z3W/Oe2DQKOyM077hcTAHOstmVcbA7FfNa6t2vIEL1v0cPStBV42rN
6OiH5ozET08gCM+Qgolclm2iOgG3mWPfbhqN8X5DrjoKUuZ6Fe5w4JpQEK+L1gCXH2AJL84dzDIS
iFzapTzvQjjCeJ6vp1uk6uLdAcHEmguQOgZLuhrngP0z72EWmtfnpGTZUnXrvc/CAduKpzmEmrAE
1Wb3YGWV68pAqj9DXFFI+606b0mokL18Ab99fu5zbmo9y9Rz0yf/BfBxTnbhnWckUoNbnUUZrn5j
nNuCyvQFqolBRtcckc2V10jUxMRK+w38RFp9VFbDnaCZs8bsrgSQRtmhyC2ARz/gTcstTeSj3INM
/oBVYf4F4M8DEooptNcoOi6h786PNCfGBeKKEGDATt6Y85F/v8jZUymbjtG8tphC1A5Jca/vrzUE
fQUY9/yuEBIKNfcMkloUpLcCY3XTk3WEDHUkaaDNp/WTyrz7MUcoGEK3BqUja/nevFBSq5owiW/N
i0neYTboqsdb1HiZq+7GSew4pghkWehePXhOq5OsSpnGTappX0wb0/uVq2O4EEDGoIyTAQz0w9/h
KY0zSRi0T3AFwrSr0jnCuh8f1oDijwnAMfe/VMsLlqMfamlkYYQYam6kr8nAN3pxmVJF7CC9GHhz
33SBbsbGEPoiaNNO+Cw1dSXeI+AKYtF1rm9ovN9HwZZKwIWlg9ITzYY4Q0ivKYG1xWBfwyeynfsm
eMQ6UJQAJ5xnOHk8OG7qxzVAnRR+TRhsFj3pJ2suaTzKDng/gUfCH4joIFaa6xWoWl+Mql8s1+FP
YpBtsVArg8QNhbV6iR1BFMPNV1bfV5Y3bK3J1pjLplduwxN0EVYT1UQtV7CLCzmSGyhk9c+OIXbn
+mDbfvpMCfAhV7DGatb9gCXiy2Hj3i6dv5jy20VQK/jmxg0AbWi5u/G1+CqBt2+xtbP2nhGr6fz/
uW5K1jglRaUafH9e0iLzdVh8yHydIKv51jrd+sIF/u+DmcM9jhiYrD3Dn1VNeeYLmWYD0iE+tXFH
BJTOS2yfHauAohXGxMjJ1dmtFaDmjqZtMI/qPgalEvHDhBz4ajpQKgJ7YFo/EtBR7kdy8dtOdJkp
RnAqM1AfJ3jdNleILCQPoafNqP87DsIXbXh80sxWcFAQDmSh28qDiFPukwbOJ6TM6xx2FZV6aplF
1sadrZ1tW5HQmwQv/AGmUvPEeNc6vhXYuPUdDIUb+6n3noq9sH828DbaseMugrhOYHhzDoBPzvTk
Yrqd7FVy2mhcE6BY0AsAlW4dKdJD3292+kdQaOctae0RKhO75HESeia3p3PC/YzbyGegnFph5Er5
e3YxwEvgjnFkY1Y3ltDRlmT0Qhvrd1zGMnUuVupWqSzm6oG8H/B2BVOYbzq0qNBKbI9Dg5FAx2CZ
ukIR/+e3lP5+St9nEtjYuZsgGgarFr3pur3OHBPy9hYnMkZsAqWoL2JL5XXQBxHk2geLqJ84YXo1
kBfKpRmRiBuGz6ZRVrFF/pIXR9rLEWeoZUSnKu1Yb+AhDilRH5mDpdTxEwd7rJ+73kxH2LU8ITed
pj83xN2MxRpPddjx7rn7HwwfQPQj+/ojnXBJQZjp34og/gAIGba8K2bKw0VyEzDf0DXMyiDBXEsJ
Rfa9sUKsBkTe8YVa40q1Yb5mhyQzGbot3TOdfXVMsOoevAe42DMD0wyMsfjKEjyYK+Cyyv4E47bh
Nh0lQnAXNcI1/aGrlKflHbVdmWux0G7IpkFs/55sgWP+Y+QJe/4ZQENqPKSVmaX3jMyTHe1QlBIw
RfPkD+Kv2QucxV7yvm7YApRQM57k1Db16D59rbdHO857grpRL2Fj+L1957J/fZRlbVT5xqrlmpRP
2vYWtVermoocHGB1Hm8e4hHZLsUTO/3R1Z3zwQRVclZGc4azPYQS4ONCYxZAminZkMiCv1ajQ8qt
J/3zTMgRBDBc41R9sVOtymo4gcGrFGRIoZJ/S2edMevcfxh/MqTnUgDGUzQMU/vO+z3xlk8/Ng9g
BhHE7zDpvE/x+LcCfPqPWGCs6pClI5pkp2B6xI6FlsxLZa5ZjQIGkGzEpvKR6pgsPSWcOFHjOdNU
iBYqVPFRdsLzuk/jmnpWdsTxf81HuPPohEmcB0bXOv60UcAKZ+ipFes+lobpaa4YkKTH8H2eQOfe
PtJ2EJUEv9xk+tAStQf7MFwJO+6bEuUl5Cs7cLNr0zuiwYvXlCCCj7SmyIsu9ozZQxC30i38Djtx
ojpX42pNvWHPJiYLZzblBSykrfj8EoLgsZbxa24V80Qbn1fIDF+AR6SqpPWfJ4o0nLhsP/9THuad
jLTkZJjdvM57owAcDknDmWpHc/9HgTuSv4jAkDgHNkZoo+uXNbjkox4HCWErja6yALSh7sOPPEY9
Cgb0CeXQGlsaEZPvXqYShea6w8994rvsPg3GuUFA0//CiKvQouwgVfOWuYQ/872AcQ4ZZN0DuUls
FoIGfGQgorWxIpm0gS15DE+3YmeRUlcHea49AUdVI0qVHnQnH/R3zliDQBHMderzL2ix+4mSjKY1
nAY0XXipwnElYJqnZipDiF7M2N2QV8AYmFGDhiWhJCK7uJrrNu47qnfXTLPsBJN/4hmecS7zDSNM
7EGfhdiuoQ8zfNJLcCdbs5VTghruJd349iciPbyUFzinYl1VVfmVAtA14nVH0z51EdZx/q0FBfB3
Rme8CN8uRNqizrWfgbzPUzaprgzKelWhDO14TGAqH6bFRNXVKzxxBVZqCGHwLeWKzCp24bRYEz6s
KylXu06CO9qQS6fyuj8Of2VbYj9p8aZYPWvQeTfMRWV2X6FLPWWCflj77Uss2VvbGpEgTrsi1L3p
BZuaICTIYw9fwm+i9I+pn8+H09HELxPqL01ESJDva3XDiXVr7YpDx2KAHGt1D0jerdUWTzRTch/o
dK9XUanimHz8+s3PoIsIPkA0eSUBzA/sehyJ0MyU1KPe6XzsbfIcnHg6QWKh5vnmQc1IgD/WgLzA
78aUxXpoOB1tr1+ebMFxUrSBRdprlRJCyLY417SxyJKaE5k+8hWvL9n+ezQinZpCdhptoFwCGd6S
IUmqQhsanPiHksIrerccViP5MnhjqXKBqOhAdl2i0iiCqanOYYJjAwxUQOFh6U6bxRw2MHhYL3it
H7aL9VRvNmek+WiEsoRvTO5gbei92rI+jCtY0pk4ZCRYvGTW+Hr6E0lW6yw+zZ1v0Ul8HQY/JdM3
gsBfV8toXhBhkMH11CjrBuKKmppHn4ix3z3ehGwqFBXQZ6+3YKgC39EEH4++eYp/dM1ajL0NrxJN
Jc7u9k3FHo/KqNxDzc4vbIrU/B0kzhwEFVKIvMNLDN9wLlQZhqwHj/qOrf5ofl23r+eUdRvmHNyJ
Ix9NMBs30bpyu9zAe0KPe6IDadQLApStDxlgAuOXR3gjvNpaEszsUB/KWo3qcEsmKW0tWEukGtnR
w5B+hz34jn3xkRF52K9HZTZarCE9hYDA1tMGqarSrYZffg1Z59n+skAVp3yAwflN31uQ79sLh0aG
+FlmiJQH8shkX0OyTyr/1WI3FBYtiHJbkFAJh0sLRCueZ/k8XKx6eumTz5P/k6QSy+PQfc1AwHa/
5URcmOVeOJzS15+VEhYiRrJhoEupMAEsWdSfDg9qjQQYV7szp2mrncMI6JOUHVQMEF39oFld3Oy0
9U9ciiAZiEhygOSXQo9WuJCdshNx0hutS3750EqcgowwDVOE0MJ9d7xQ7+Vbkzo+WhcCdHKCZ8xf
2VwBAZnsIzicRXN8fcOhAs78r976n945EA2aKRAcR8LA0osTTi8U6uKbUeHIc8yLZNgITfQmiQR7
9t7a0ste4RxLvHV645u8YhTs93ziNqepcADWVodgccP60+k3e/dbhEB2i9tp3uxLKvdrYOgOQBuN
RwyShejH1SR8CAi+03HP99zxuLacyElm/Dbt7CeXf/aXpgSYglbfNeGvPTVXnTqDrM9L/ZJQed2A
ocPA+Onha68p5wmZCcooUEosYlSDSbm/D15ORgduYurTg/h/rLQSgstYkgnUdCVa+3SRbIJTisn1
THcurkRrMJxxiM/Yc+14OeT6HxF2x3IX70Rr9enLN8DKrluPceQ3/EyIIB1cyeozQvxDHzK8dx8d
4yUTg4vRrA1r9kdHm0DnZ/zbBYXDlvAabYHNAhpoPQrAiakhEMbInjYGevTThnC3XaA2kXBDxUO4
q/ZxN8vRW3lPiEhIOBZJe2znaiHQML2BKp39JRLeLRzwoCWiZlf6z12pbYqxHlDTKT4z36j/YUUA
JZ5iT/HiO6EAC21UltIw/KHuXYwiTe1P8jNHlheMeAZahK7N1TJBY8XLpUyyQxnoVtQ/kqneb/+i
8uAxH8uDlzNQ4XkiD647i3/KhOZ7QXmUtxA2RumTofP8gjGuPg8OJtKq5XwNftuxJAO2Y+6VCOwJ
8mIZ+vC2kdRi/hTFjOMImQo/f1+1okRcfn51a9X6jB4gQBZOdyEf1U9F0gdSaCPBu88UxGyRL277
zP5NH86bvnO20vakIifnBna2tGQGwOyOYw07kIyeLJC6B/weR3dsiSmXon9DVHK+yXt9Ngtksrq3
xvPfzNrK+YRzxixWsOxGARNH5zibP3dTXvA5GyImVFK5FIqTSkX9EjiZz/VlCEESudKeswpVthoe
feFWYjYxH2fXWrzMl5ZJ5HKIi7s7AQlnP8gXvBL22WJuooth/ttYU0hUb5TNxzvfPwvYS+oUOAXt
ux2655TYl/VGPMcUMo6kcEYUSowIVhvl9gI749tpWpPpxv/4vm5U4lNTEcQcKFpfJU0fKF5ao3uu
mAdZg6b8KRUjLUydK+GCfOG19QQ5gnq5NWYYoGFQS4tkQM4EemhAd1uGlWKX06oOLRoZBTXYBglX
g6JfNAl6rl3RV8Y6vwBquKQYR+Lqzuo2WDOAURrf6eXf4zVcw6q3bkQpSbP2KBQkrgL6qQvjabNI
KKD3FfD0GcVpC3Qp5iH6n/4cXmfAXUakTd69s8AL7fksm1hWgJ1uQLwjYDmbmyUnkSNHJlFgmQg6
LjM+JnPrO+ZGUst9rF+HZ2aiWnM4uWESlg3eHLzNer4Qm5YFd6aRBi8MUphPxVt5jxFpUMImsiHR
uPStQsW20rctYxEqtQCEY2VL81ML3yUkbvi4nVlNTMAdeyx39QQJDRkZkfVePVbFgwrfJipNWHIQ
AH9l4ZBi9VEDU022340fBLsim7wWT8o18+N2RcwZVUyOWd1Es5KGS0ZVsldIx1+yT+5zbsYj1clL
JaCJR472ZC0g/R7fyzydzc5zo4X29lqf6TZSMlmw4JEAfeGJ9t8cqdGJ+0llusukSpbZMdy93gUX
rrSE+06h0u14U6TKSE+NtM2DK62++qq8vm5PP0FahIYzFF0CVwkUInXDUILHLB9+QLG2EZCWlPa0
RoZcJ4J3UUMXfVvCPC5muLPE4h2B8o0deYeQGw71g3s8MkypQxgbzqmUvKbpwRiEZFgn5KDKjmpW
Bxh6/pcNSX2yRoUp/loQEUVns6YPO9gJSDBHAuxuw5zlPqbZSYBQeOoLf1cAEyzQnCO3VaGViZNK
2MKjs079pgI+OMHrsV5PzazPliHtWO8MHXVO2sOJGbVHfb0h47HcdkZOdNtC/3noWNrOJZIhD6pW
Y8zdriul60yjqrrpxRoLcJrXA+7JR87VLBYwgH3uE00Y577C12eiENOl0q/XeLxp0YH5RtgxzoAs
WLysiRmRWDzk9J/F3AoLDgODm6L0zsn9l4Kibbb5vE+/Yvr6dLX/QFIkxyRzp4gQXuDRdw1qjTY8
xNA0C4wAh9Hf++QNgm9a7JJlC6gUNKN61EQNKRrx5X9k7p68yizOcRXNGwrjwiHw7EkcpxJ8I6lj
L/junJYm4aZN0zEqm+YcNcV7Wc9xUR/y8cb1y8BaMkCjf1XiQAOHyFLSGtbamyyObAAFrdIXOxaB
3rqdq31YxSePYRzKjP5JFuGBiU4Ds67m2DZCPcJTT65dKdyZJ1GZmi94KdqtxP6oWiB+luOUZ8Zi
on9JDH4qx2llFy4p17D4i/o5APcu06HxXyK5oTQWgPzlyRwhTNYFO1hp9cOviwTeCg4SD5bPPRjN
UL3Iusc6dB45YYKq5NzKr2QArfsq5pIpnhrrGYOJI12hOrNVmyWJUYLdt5XN0bLRNs0OPqyijFBz
h8tX+4Sf82dTLi470CJcXTrn2HSuk+ABYsKQKTHuyF2s/naZFOOkJanyXN9Fj+q+4pyxVu63AfHE
1QkxOl3U4rUsOPATuwF+uey6RiPC2X8VWaRE0j9ZlwD0C76Uh4OyymY+eFk6xPJVcbBrjlzI6fy5
pM84wWRa6LTB5RQ9tOJtievS6xb0VZQH17Xu9VxGXoSem+ai554Apz0ollvmN2LCSCTD6ajsBQZn
Dh8Z4Z73mpMUG2JvzZDB569RWKAOFixx4Rj5kPDhsUZqBBjToShz2kTxigTDJ0QI11sIwwWZ85Jk
+/UMhLVKK2MkFAtMIynodPT+RUq9z7rfNE/vVfGq78eaCB3igEuztkaCw1AirSv51LLRPoFsrgHy
wAhHph7/uEiMvKUhpuRH8fK3Cr0OeSOlSVFwOLqxTJ2y0ZzCknHy4BiX1FLxO9ubx36DLFEZuPs0
5PmuDz35pWCWbEr40ZgzTVeUFRc2BaYIZ9CI15zatmzZa/rgIC4BagLr0AuibmVMeJ36ges6fWmG
3w3z4j4rj8PFq29jPaEQ4lDU4ogFCczyoFqzgwfoZXVbQ7lv+wW/3Xn17hXTsvf1bjTFdEvt/Rpx
82FSxkva/7EL581IW/6fnhoMCPor54lDhasG2AqyyCR41ohkYzBDH8qG609ASF4bUTAyyzKfkkQq
qxUbxt0LQxT0jgtcH9+3uH+6mBwozKfw66cDbTBcKdzf2QBbNoLmoMrKIhqsr0hCLGtb21djyxOY
DtSjJQ8exrQNgCpAQPNwi7LdOhYHT+xQGud8wuKd18XYtt3R00VWB3CLF0YEOZvnDbdACe0z+tGM
4iILwkcAR+hiiYwLcLGOjYGAHoIjyq9vbbFej6/8cT1AygWVVA6Gh+bmIyUCIEd0hwDJjZD7I7k+
sux1b36ZcK/uV7LO5cQhWz45EwAv/UFv+zquudjYvewSGqmSAQZh3Lrw4Ns0eKe1iHBvbfU+c8wD
WQ4kQjKfT0Po9JNZndibPLikxZDEwC+0Kkz/zYosQxwdh8tqVA85iSxwPVGOXJDw1oje2KlYilIQ
2yum5VWcwbKI/Nk1x0dcXXKiEPMXpUPlr8bJJRybpbpjJ9TPRbutWtgi7MdEsAJ00x+zk2EgmEcB
sMmFQkEgitsc7zCt6Uc4PI8NQkQvijSDE7EZcRU+w1xVtfWg/uCR2QVcfaAeA3Tp4q/Z+7VTI1lK
CM8XQeSxDjTaU870kyH/J8fhZ5LAJDps5kv42FVh9hdyvlvrG+iDx3emTbe/xRbrb9ivnOX9er1X
xsUz2UDpFkfiHhyG7ru9p4ZUalJpLpsqoRhP3WepWoekK7Z8fwHsFY6322GTpq8ysOsRd5S7dn74
aDbkX3bnxdrdVQpcgkX2UdfgG1shwRY9h71MDoi2uHDUvC0Yz8NM6aRyrcRI/hLAmlfmKVX/zNJw
FgSldP2FaMaYxgekNFIHCSBW+J+jR3tXOR5sFIKF9ny7CjT1V47S7pJOc6AVIkOPwQYJojvbJluh
2iHqvg9/Mb7WNTvLq2u8IjTHXIw+JeXXlfGFbnCylKPKIC0PPVUBlV7Ub7do+hzszzGruzhyHPdJ
LkgmL5VcCvWPTgrmlcMjMEhYLOWRh4asm377zTX/0KjGGx1OVZoGZVzrpjksANT3N0+hS+WelVew
T0UOJLGFDahLDYQbiZrHzE1xpMKCl9TAjCWjDxiTKYXqI2v7mV2KJOYJUWiFyJm84TmNOpJZ2zSi
GhgVKUN6YRpFitKmRf3YFERQfNaUen1MmgXd0m8JMjPbcfTEErW7bZyP0eSso+HqaYoZEh+YNAPL
AdnoVh9RRcDJgQlPIL7LPRjgppAhreY1kahyBV7r0l3COq2iGeAY6bl5IjJwJQpLJyNpVXXyrlkn
YL3vncw9WEtxjcyS+pUQVVrNu/yuJP3eywdbd6g/tZGUXGYs/ox+eTNT3AZ8Anooio4Qyr43FU0k
A4B39LZj1XfD16pssFtgEpakOKvDQKsfqTvtSNBda0E8ce97uc0bM7SXouw4u/9UFUPZ9cytTIR5
TxeApGe5o7ktVrO9kpXqVsCk1dYIa6sA1yZk+A0mjEoUyeGse0/zd2xgwLJWlD7ZOU8c7ZPPW/t6
MG2/+eP5Z2wWMdd4yRlpB6apf02eEcDAxVfyZiDY3TeDQkpG8Awxh+W96m33fyVlmEi3KBmLLyte
VqgYbnJWf+Ovo2jSy+OoxOf5K9WFFSVAlqNckHOioioBgU05VYzWvpDN4UaQ73dvVdDmrokoLNii
mLNzq0VBecum2irb84rD7RQtmHt1DP44LNF57oW/Q/N78CKIQ9tIR3jEFbwu5kSBox/qPX4UkAJJ
sew8wUCs21ECjJHjCPBLz5niNPMLsfkRD8TonWve9q04CiMHRZWKp3kIMC0OVj446gwu/wobvQvo
DcH1MJhMa0XGRor/xhSEGNTs/J7FocSbQVSzacdPZkoly+s2+osSgfxTKagl9PATqq45LJHmbWYm
kPddy73l9okxCdf4la1xcx2rXTAY3CLWSZD4d8iZndfUrlVSz1MWM0rQXniPGchJ6n0F6Afot6hu
w+WSTLaMRlNd4LV6AcJo2x1GLA6HuSoCgfkR5bj1Ufam5n9dM7yMovf4x+8REbOLndTtRP2CTxwc
leseymnQY0CA+AnU4ZjmmHrLq3EI9oFDhUwuvrptKEd7MPPUDzh+kM5xeDI7tNYAJoHs2SS5+Viw
qBRU1hk3vKJjHTuss/EYaz8RaATE4fXWW2ctVQ6xg/64lhnYtInDMbfz2G1PDkS7Ib5Wf02SpKO4
YJeL1fHWKKUYFwNwJ/Y5Ad9oSd5vfsHNOrEBVIhHlTRsE1r+MtCzmyNXGscaNpt9uSQWM5ZqqMcv
azeJcWBBm6DA5MYr/zH3S5rpeiYzsEJ7HuwyXzfzYVBlUilWOncGMz5UQTe01F+ZfAJeMrtiQYr4
byeYr1XpASJ/o4t9HUP9rRL64tJ0PzYUHPaSA878adFi1PIgo00ptjCRAfHiIVW3QlIYFrCULQij
0X7msdyW4bojsWzUAi+tsGgnkr0LVRUQHv1FnkZs1AseobGNWKlnrbX6Mt6vz8jMk/jBjSsadV60
k4hQFawQR1y1KJ/+RSstljMqeznAcVlMUATBfpNMpl1K59+ol6RqI1ojVA4TqSo4CeF0UY4mAXhK
D45dNSQ6E8gKVZgRexVN27gIP0/qSdYw2zVWnYgA8U6TmVX9Rl8HwhOo0MGiQ06MT3jOtPprAO/e
egweFMe96c1PxUapLHuaOLYi0hExnYLpM4Mwl7vB54lDQiGclihSu1SwcAku+n+0R+ezZL3E6QXF
Sj+DP91DBJR8/m4Ng3K3vW++hHC2wLdv1R6BT0Q4Ded+H7RkRMEuFOEDtQTR8PmHIcXIe9Pgc/+/
anLviT0bKsThsj8OhFPgv21jPbCo+QiSwp4tlqHVtzgsS2BwrTy43uLZ5DIFa//pIfcgycDP2Pya
z2Pgnrkujg5Q0YamBnoClGYy86JbcaOuBF/6BdBw0krDNFFftf1oXGTRdhDHrIE4b5g9TrCE31QT
9oaSQE2OQuYzDvHx3QsmhLYL/9hgZdSLdQIyZQhwyMR6yYDsoHfcIX+ulpg7zN3djL6XZTHMdljy
odmoLvbysmcPCZCbd6hXxQBb0AxjJgSohj/QbhJWfQapwSMJXfTmUp9y3dW33OuGKZ/PWcmB9g5G
zi6IM2NWelmzq46j2z2KZ5TON+xoyNaLKDJBaIRdIBe7fZVMH87UG8vhfSASnOMT1nbupWSzUWsN
AK6kcWotI7YHgmfMK5T50VqpEdZ5CFNZr2ygUjNf5hcca7PKQ7EIIh00AYkJLP1c/pOL4dk3oCd+
tFHr0hqSnYEGcrbSBUuJDoQWQXWP0IDpm7M+daF2W8pt64Kf8iH9CIEkXk/7o2UAiN1P6/sy6jJv
awU014+3GYV0bqvkEuQLAsp+lJP0JpD/yJTTowDZv1qJzaouPUDQW5OtgAgWI1eehuFFITPMhU4e
J7cK+962dzuT4efeZ2EonnoOr920t3Es9gZEQt93MXT7ToQw/zKE8FTuESnnjy9/QY7te2q/1uga
HcNUZySbZftVtAUu2QOf1tZbe+cKlreSeGaojuLjZQMSthkFqQB+1tXDX9rcWCGsrhDa0MkQ+bbl
NnvXwdKtUIyPHMXNfIpClYEjtj5eAorJJHcFNApnHglyG5UZODSfWgPH1oxzX72qkevqVKaQhapT
2J2zQXehtrdsqa6Ee9EzCLsEdw+kzl4UIdovOM375ahuXigacD1v6Rv0TCni83rOf6Yltq+KMKRQ
i9eggevEmPqvTsxUGUpl+WK5BDWrbNh+6dmOzZeVmpO6u1oSevkTzeOrw8tY6gnCSHjGn2FrOwlS
a0aSiQS/0V5/6Ddec/gJc52YsMrj1j0VLePmcXTSd/QQMS1He/8fcXM0opTL+nC19f5W/G5XMyec
x9oTzw+D7Exs6KSrURMEuH+hmmEaBT4UPvrcTC4xWpTlT2tNKr2eBmLGYkRqyeJ23N8tXj5TJ7Yv
h/ehQUAx8ml8MziXHVmEuECCFGBZBuByhTyc1vZ0rYiFYAvgsIKLVjgzaYNa+ZFzOB2+rIaIxo2M
k3qECkYqgpGUSJtTDSlzxuNYqz1WGeNMFBTN2t/J8pCcz/Z/K6WDXFZtdie4IIle5KGqQdmmrmB3
JcNCAdk+aIZDpxLgY/vOqR0YK97dk3OIjGCrKoZbtQPzqUKreVMkCaa0A5FnUvMX8UquXtI+y8Kg
2ffisSejILNGTHrRIO/U0nU7ZnDqhFf7XhRok4xfwndIm3btS+NqFAh0KU44wvFAHhAVIVXdf/60
ZAwSQwEMtpII5PTex1vy0+aV3gvnIvlRvDaT1hMfX/qZ6WRJwNQVA0i+sBSONPOwS3ZX4scK1lon
yJ/IvR3TckmBVLt0I5ztKb8PeaIfiddQdcleP4fDNdyxxEugIHdC4U2pz2vV5uwrAlqpSIL/ygbY
985UkVXNqkJITNjamTcoP45jDjE5+nN+psNsSdPHjLMluzYab8+NMMpatjPZa+qxTSQLGvkOufU4
fktJQDKSa39KcE+xG6nbqsMaUBpC5zLXjWkYQjdw0xdv6wd9u0nW0u+rz3F4BiLOxTwWejMnuz/i
wOD3SoovGEgO2R9HU2uw1lz8X+4IbBIxt1ihUyCo3fLkVW49QrojMQ7lrEGxkLIOWzWQGe8uWlYP
Acizs62Nf0qlqPmKBW77gIC4RVlhFvO1eplv6BBzS2uwkELpabwQ7g3j0NMWdyr5CH7i4n2LpaeN
Hrux1xXjoZRLyDANV8ytQIkUKzGxV/gKqx9yhf5td4wfPPWGYnpoJSCi+ZpR00yywcWZ080pfl0l
rgkLKUmbFze6n/08/gkw6eIitTagdyUUJHSiA9IHREpaS3flSe62nHxox4Nhw9mGK04h/jHVgq4v
SUeafwHErD9ZSje/S6wiqD3uB2Vg/AVTsng77OODTWhC30HRunR7Xaff0SL53T4yG7YVIWdUvWjJ
2VGutGbQ3L8wgWefdV3N1eWPbkcHEKVvXoHpT8CCrbL4uhLZ0JFgnNvJU5RIhrNYzlQvBlxhiXLM
Tb4MUDn//2ls+QUOgM6yNdRX3F7n14XZJN5Tkw32YdvQBdpKgB6F+Dvu5KR0GKHk9AnxevgvGNTt
XPXGnW+tE/0l41q8lO8+NTHvgh5+896ztojFEe4okiDVjHgWacgXOt8yVm8cW1mRAYxD02ftDZlQ
7fNJje7UYaklYMpZXYqq4hoY53X4zXuU2wTyqEf3inURqZB2Sdr6Yp8e2XYSaBUo9JTXYBAXfzVk
1mzZmLV/UPND8/W/0ckbKRqqqGxKTP2pOYDBIh6YF5mYwB1Xzl8x3VSzPRgKxRblCUvR+nmc440B
CL+2NrGcEt2RdJhfYRZ1w6eZGE5a2xtjivqJnSYM392mWdF6T7jwjgESY2wTyKcfb0YEvN/c8Apx
AYahKvkV2r2lVDJ1bCI5rrZKxvFIjBJN9gPDt5KQ6ZO34G4PmdKTqTzT+28999b1mmCDhO114XMD
ZkZeDvgOiCxca53AJzv2xl1vi1bzhcK14kCYdAlFN5cPJU4qknhRbJR55LutknffCeNpJQH03G6Q
v9wTTlNDVWwqc/kDebFkwxmIo3eMpizzS7pQeExEKwXKcvkKTCwKNWElgQ5ttdLqWasSd5PMcNq3
xn3dMTMB3tgm48p/p7nIvQdluo0yZZ4X8Uzu5HOP7ANyPT3y1ZFGw61ThkfOBmf4RfploczkPzvZ
oTVEKSeW5UHKhB8fKBBZ+2Zx1EyhFm2SdyMUfbW2QAvJAzhKnS2ueYc+XJoahe6K47ChEzHTVl7p
bCi+hx0S95+XbvrAQcvStRQOqgxNf0/iKKzAc5X77TmVVdFgi8THCfyYSqkCfAyQ15JtZof1qNjA
MahrfnCstCG0y5jBE6LcrIuIg3pIMh6iE0Bwk5hhClfv0jUGTCSX1EUJuclq2zqNe8n1BT27SNEZ
oZqg+WWxr5Vp+tn2twSr+JyUnZr5MjYCxe4+kXK+BBOzqc8wUzvlXwhn0pkmB6bUyQPv9ZXHGt+q
QMqyUpo1D4Jxozv+Hf9ZOpAZupojv99/zTO3+3XenanfZ+2JLo2rKU9cqnatgtJIjZUFozGcscmY
0BruvuRQSOCQaKEwJTW+feoFCreU3jpr2X4Yep9I78xKWB2hJqkbOrBuQ5y8Syzv4jGWJXRYAZl+
JE5Ezu1CmXxHbVDaWLAaDXf3kb0a2ie6Wb7eUFaVK/uqyuRsm63ECvQiWobxGF4ncMAUfMuq2V/x
Z1i3OXWcsBiqVPuVZ6cmvQC0rD7gPJfJi2KH27nneseYzTaRupqQ361uUBW8zj2YjosvQFyK6EgT
Eb+yO8LDuifsJ/qbPWAbGPNaGrK8xMkXadDIwNfUC+if+ThkrTBoYESWHveGZFFgJxEErJsf4xyy
041lXACUTtcJI6Y0nCrZv1KV4CNupx6Y0JKrHjEhy36eqOsx6ruW4DJhU/vQUZjWEVl0nGfdJSJP
NaBqTcezwBBygDqk5glS/+6SpGUbD42J+TXwW0JNAOn0/8JnYhmt2GXbPvjw97sBgrbVsSMGJoR3
IU8KO+kFfo8tyfQXr+YaowTlIN3a+yaXac7ZcYZsJ9AodTdkQ61MQOcKzCnvd26eRivzN9cfEOFm
aY6+EHs9XCFwKKT4GHNOxTcfXnielWgkrGUtWyRNvQW923z0ku2/udGd6Ovp86p15At699WyOrPU
b9aFv8WacfJaKjhQGZgclkVxC310jb+nXinsl5QXmB7SLpapUQGHUz6W7cGgHE2BL1Xijwsl4zTG
9jHcBOP4jYLTzRevr5emlWV7clzzezU3aac1sexsGhFfpBjJ51ZDUjQOVtr9J1xOwY5GJN8qwgUG
Gu10pzfaCBPNfaofT5Xnfs06FBFpHxLVXmKsoo/eNvL2xmsTzttnvGrQdLACTmH6y91sA+Fss2k1
JAa3y1lNMFT+91mWwCIIUpqbWoG3EtVwDy2tmIs/JS/xt6gtPIOE7cLcdEr/j/O6FuU81hyFLtpu
LxdjOoPBXdD0kCbupSS6EBhZCgW9tCS7DFj9z5D2b0B5sNZOce6wVbI4iy2SqkN9KfQnMuR8pVt0
0g6Zth5s2vPdQWkhTG5gKCtB0eYCbth9Z4XWy8gDS8ewNBN+4aibijnIXzdCzbmd4stMga7S625k
pXetpcjnkeV3NxKKv+ChbXTSmUG1JtndMS7iFOWCErhvMqrtlnTDvM4LJmXGeNfP0u0MZT5FyZl4
grViACQZaWk8kTmN+lMWXusI02NPRCXrtxW6cEqk4XKkF5mW46a3Zmt3LN2VZb/HRT3C1DEkG0Nu
FVkLZnkh7QAwaqN09wgPe5wcdEtz7TeOzuKSYhfLGL7BZJfz9JxNFCq/aSlfGnfz1y89GLhCDRUn
ogTMoLb9/59fGQLIaPlIKR13L5JlpgYiryQpvBxq+myoxx6ET9nLpeQa/92v8+T0ztA40MudTvMK
F+HSYXF+832QUFw54MuY3BEMhN7jxbzlJF/ulhdBRJ6ibiCb2O7UEppD2lZ/uZoU9YzXvlWzx4FD
RPIyjOLswewMtaJwukfoShYa8EKr0zBekBrSVKusTSDp2+Y2NiyG45lpuLfglWnUpLeIQEsTvztX
2zHeeoUFZ0tvEmeSyDmuibiY6U3NPwWr714wHpQCCB3BxaDXflg0fzaN1Y5JQ63s6z7RPftcwmDS
dbpUioLkzg394o1gbVMeqy7b/BxX6CFaPiLgTr/YGoTBjaZAX53gvK+3f3ox0KrZrOwWZQ9/58L5
uze11N7qpscgLR8MmKWakA5JmFfDLO+TZ34Mtiasuf1r2slVOXURNf/v4vzTz3AmEOkVyBw51QIf
gnxZq0KsV15G0niM+fFWEYaBYuKCdfGZhwOeMTVshsI2zMItRxwsCD6SjulfSoIO3EzZXAgM0Rsf
ElUNBggHuj1iTKBBPuO5xDUZQJunMwT1uMqJlIzXBq/s0iiO/SGjwEm406GVxtCG5PNNhxN3CwcH
dof0AmNS2/Mt4+0MsomY7UK/07SdNiUb796hu4bspkiV/ZpaMpsm3nrofLkPoTHlaLHPeBuDsF4P
tIjYQyQVdKqMYKV72V2/VujTX1CBaIJwasZyu8PGzB2aXudhi33H3QMf587Of1SI3JO2caTMYlSn
oKxCkC+CiLArEZYlb5UMgP0BtTNK4PDpbl7ZqW+PDvc2nzPuHX0MJdx1HMbLNQt3jZBltexM75E+
xWx8vXYEeyjyA03mBAUW5069YU/jggAKe5cvmdu9cKp4pl1EeGrZmCtxs3xdQU7L0iSUJY4auEQ1
xOaolrd1pFEPSLUBzAErx2xUkvD1OT8BSsExPod4p8BcWVXN73P/gPb9S6kHwxJEEjusve0RM2Fj
2tcsYOCPg+QSfUZq/URaT6Fb6rcGXLCSZ62PVpnN44Yhc/u/vTYFYLtDS9B027+e/bqyIuKzO5XS
1HGNTQPPIr6foknoii1H9Ftk05BLeu4wv3IU9gmCt388tGLQQg5379Cw6X73KQMXsY97d5Zugu0P
0c9wNBmlg3shGAhEnpA1DYuNe1Vobug9rTzHkaSblddWUE6uqmvZUPVWoISJfNuH3DJqei7XLIhb
XQuUwVLtgqphN6gRnNKHKyUiKZLZ0zLdEVALG/7YDrpHmuwOdQWLNfyHFC6KVDPJQS7t91Ef3kbO
eD0X7eAPGRTSCZNAZvCpTDaU8ZhgRDRgmRec/wx7tgFT1IzInql+O/25wFJaOsjMAtbJK9emDt/u
vs2E2Geyd3EdjttVTtTLDibPTmTskoOmSdRL73yz9h4M356k5pnZpfdFA5y3BkneOGF4ncmv7fc5
QQe/S92dnmWBNwOz0odhwxOSvJcMe2SWm5b5bE/Twic2QaudjvJvYSpORQPighIsM/6kvn7uus2u
347fmYqE+4+a43mXpfDTK2+WN4Fk3625Mvuc4n1OKo8EnfqOkZVcVXd81VsUV3rJq2b4tBMtPBJ2
JnOfDVeLY1nYpV6vuKfnSuA7NOiX3KoprII/IQA6j01UMrF43L+Fx6x1gXxsjYOn9bekWFb/cp8p
V1i6QxSQPwOD2deNQZHShlMTtzgCdl+A0sGLuHCLjSBNv6DWHr1+N9xEBGrDDAgfvKeGtQo+ZWJI
X2dKbG5XyIICcMHK0QDUWYsMNeTi+1vTNoxkoPwDiL2N+REBA/P4BNYY4a7tB1/lG9Zcllc/5h7c
C+P1chnzokC0ZsuBVHLPHOrMW87wJaCiNKUMhFdby3lWtrspmXllYEORotdeJnQbUHSRNUUID4UJ
pCSvW0rN8CQSjQYCeGZsaKLxNBRfHoyMvli7XxMFmJG/49NNhZ/X/NUbKEnGhH1WyyFmcU++aYY7
ezD6E4doLDjX1LJUi3UxJ5kQkyojrm4M1KGwlL3a2oSv0sYOjRkhXQtRS4jpNlXcN1bXBHe5p0yW
KfEsxbF8zxFC/dwMpUL1nD7Bq0wY1PQJhwOW8EeNKaM4rBaEPFG6ntGkFQB8FrJIK4qmS3Pc40ks
nwVFb5kZoeoNAk1+K2y2W0UlUJHjIBhWnqIeA8i8LvUc0KTP2rSgCJiz4hLdodHiGGrci3G45V14
NvrgzKBX78l2dwgpWu02QA7UncLsRgznZDTqzhknwZSDcAcY0n2qA14O6yFTWFbcBv/UZPR5leYi
4hNFllvD9Nx85fhewHBcuSerP7ZOME2HCUa/HLqELu/G4q23eJd+RVeWz1BbFhN9OFcrWqoVWDqK
7TrrC5yC0jFQU6eFg5ZdtiNZV6XiNsgYILhyY8gQdelCRHHxVB4ZCewokTEWu+S49R2JOywJxgSD
3WSPUYYng8+qxtwl2kapw2FerdTPrWyBtg8t8xB8ZVWX4oH3hMsxRVQ/dodDJoE0/CinHw5rJn/o
u4q+M4mU4c0mgwxjO2r907iz4I/OcxaPproGKutEyaPyWAXR71wkZ7Jc1oIJHgWYyjt2EENUo40/
UdLmvdW5yiw/Ax62rxLrpFBC+dUOZO2s31wgbJptrsN3pDY6dibSVtq70FIvGV0xoofydV78Pur6
qMfsnghjdnek8JFLOAB9Ra/QCvYF6UQ+T5L7UYp2P9mnWEAxu4o4M+22x0j6LaCuRq5NYFODpWrE
/MczCz2TaKhkdSj/P7Xafby3cCXTHJ8I1a8CaCB45NtqkdJU7vVc4HAY+vrMk6xygoXRczZAWKqp
WWUgyvTGNiFqLH8bOI/VKdMcpL4GcgBQPen9brJ/nM54iVWODv5Jc3ekRTWZlQYQI/Ke22lxZ4oq
gRB3FtxKpNBdV4ihNxxDeQL99fpGv924rqGQRdOslybSoql4e52gM/3YaoKiejQ9eLMp7wr/mwQS
U2BZwMeva4+zAjQVCI9QezV9Aym2nZ2oUY2OBLov4G0jhYGpMbyvCRwRLK1mrXXXQxBV+8CeB6r6
DR3kXhGkDIw3oRSjpxsYxXCll8sCq4+Do/LmPyoHcbBE9ABOFcvWxotjJozmmlUR6V6aCw+Vdssc
xPW93N36tOxzXSxJ7j4a2iiOkUfu9MoJbFZr3bnEvDvmtg8+JjpSTFdVcp0qJSforuYEs9d+vCXK
ZH6HEeOlVmvnVrSi1m5B5wk9gdbM2UYLRfQBFLCL7D+nYvZmY49IXYTrDb0MLGc4gVVuqeJhWXON
9dPrXxgAxwEWoNPq2mC7J83NKMPVfCCEyQfqJ+JkPmcC9SnTnE6RuQmQ9ZIXH8EBOWy7+kotWUBl
7L+wNQqgFltfs0bD7ESUNyG9t3upigUHtxDytT8EYPbpkDJ2rianEJtpq+0v2ig8kQmecmyzbI8O
QMNlOwSOyLcIe/Bwgy5lF1twJFcBlJY9j2x/zKCJay438Cdy6f3LpYgsj5K9Q0i34Zfhn2V71Vv8
XldYRDevQqXjwQ02G7uLlkuiXmJJY0a5DQJ+bT3jySNnxLDgz2y+pRtGh9LD6kDfM50tMBCifpX9
NgSL0szS2mxKPQP5KQpt4cs6U7L+hUeabyjTkQwabiPntjZtW25d5nXMEp7Q3RfmcW53oWYBcmv2
hMjSR8s7N9AhWaR2N8wK9Kie9El9hJtj8WHCJ7YjnI5UB/GtnKVNvp/IKkUTvZC5rCjs6haunGK2
lFHOZKTWzKT02K59TAjo8LYhoa2CBZLCJkau/MGeFc3HFOQGp92kv1Bi5Ypypf6UeGpUCSaHmflV
Z/OWzFCmjI+vOtV5Hsfo8l9fspwZxN8Hwpr2dsZld83Hyk37zyHzpxwqlniVudhuWGRtA+EZsNxg
wt7F+6gDFDkTaD4swLSQz7vAwfAYXoNdze213umg6HTEyBQX3Qp28F78Ha04IIV3l2gX+xkSZ8zu
T7Ag6TT4OTgivlHQvpYJzPYqnKYOf7rgzZoka2N7jyqEwfd8nOQhEX28yZ67qBzIZuvFGyAgyBvC
Ir474KIlO1X55K4wOvmldMtpMTuJ970guVAbh0ZC4u4eG5DsWhBKtxMsCVdpHdj3gVcS/D0S1a/k
DBgb5N+8uEvlYDP7cwXvNgUZlzzcOZipEGfk8F//WNmjDLEZ7ywO3jMxR2rB+nnhiA97wh4bOz3o
RuZyDWByB+1WIMmSm4rMDJYlvHWQx8ZzlVqPALlm7n/NzupvX0X98EFG6e7bjn7VTcIAufwEW1YF
DMUMpU/Dj5p4putYhEsdHxxH4a6b+9ji7GWDJ97jrRy+t1rFDmiZj0XHhSlBFnhO6e3BuR1qzZJY
CiB3UAwyNQC3TpjV3xzlP3XXAEJCvdkLyJK+2K8jagv4jXsA2EXbJQog+b7QEFc0wcvgS0vz8Rzq
A3CypSpEF+XY9qLWb2iSVikvjnXLZwNf78O9G78cLTih9qV+kYgZn5EF7gQMMMOHt7XYR+J0KEdn
Sbd3F0sglCUmhIWjmVthDWARLXnid4E4hZKCo2VvMZ3ucNrIHaDfOZMC74yf9yub4/c2E+zhdcvC
EmoTulm0cmjtX0cUcJRBuN7iDvx2SprF34TEMe17DXaJeg6HDglqATvbgr1pp3BS49V+Jm2M/iqf
463xA4KENZ1VFTuH+apGCG+CU52Bmx/yKBCpx9ljQ7ru05qYkM+gu7EMUR4G0aOUH/vozZmzn+ai
52JjMbAOh1GmuA+5sdxFbcmY0CZJzb1LNtwtrzck1pY6jRzLa1K8ERU6HNFJ1xy36QoubUA2iVcH
fihGF8zjmTg3+Pfaz5nwREVvivKOm3+DZMUZ9yNF8Dp20fvJzxLVKVsJF6Y7R46KKQMjiC9+jM3D
R+LRqUbwWBQRwI7gLI7lalC/pfC5xUU9CcLqr5XZXQ5hUNDyBl8RyRgoLuts7KP8YwwaBcCUGwjv
MylwAG50u1s886a+U8Bm1soop4PJpZJH7pMPQCrfLsFSvTfwFIMmQQULzPjhRWpitokTnCx0XDAT
fAJE+PdDjhnU7SMJ1Vl7C+S2EujZFQRCuOtCiZVnoGFaZJIgPOMs2hhYO7MavJ0ItGT/dYGdWY4A
76/rpWr12Ifgy0Y3Qp5ty7NYSose2zwyMbjTr43iwPlzo0g8ukpMLhTm94WlZLjF3bwYesvNhMYg
wL4kykm4NZ1/2tTnO8MnDXsHBd2JOBbiTWUdZUeIXmwfdK7JUaMxK9Ok4rD6G1bx3NnZbII9s+un
TMYDj2BMbCfSGP9Q7ZO5sa7C0ChnZZtgJC5bk6ydBCmw8EDxqpG6Kqn41tF0AvrvsTB2em89jzWe
325jIr81njpLDx7+4FNMsejqUuDQWa+JTUJ6y4DXZd3PUICgSjpAq8kkMaSdFEx7arzzLfPd4bW7
XksBye4AbSo2M2sqQl2FhPzrU4FqrzLnIudX8bcTBz83TwnH5osS6gaIMXuRrDNd7a52U2lzU1XD
ciuV34UYfXfRuCn7LRrUiwU1pkJ0LYvVfx8luTb+Ui9uxZZJjjJB7SnDNgkcU5aL9h5fI6mC38nO
6B4xMgyJ/wMbgcM2gaNSKp5Lm6JoS96+0O666uCnLkx50x/ENYRv30U43aMCaJkhy2k/LXJ1eh0o
PkiuV0qhcIqiHsQTwRX/zDBdLDhfyRpZ1MeaTpvy95+JNlY3yXVITsnGfuQwl43P3KF3GYOs9Ah2
qz5dLkJC3YFKPzKucTDo1qPmyTYQIGMIuvxesR/DzBmhJVvdR1Se44jN7C2z9WnLjj8RJK+b66rm
FVdw/6sGbiHNi3pnim9yWu00BUScij6s80w59K2aPXpGhqG8iAyKNqdWNCK0xIImBgQZCImb3lbB
qHpJZL4PGqqNWt1DVKFdx1xmYITWJ+UJHefnzSpReCh1wEl00qrF+WopyPU9pycSL/70EqlmzhSm
O/sMUn3LqzwSed6Y75+6BkDye41D4+9iJQhPobKUuGHGiUJdQywbsdsEN64Hc9B4TTTPVydl/ZP0
EGgFaRXxwpfJaHY8E6lsRygBKawIwtk+AojsGfmTwlA/b1I6Dot4qQsonwpAUCoPQlIzSlo8nPZN
10EvSaTNhUlizOmC2vfrDQoioHK7ihEw0bq7FWBukHqVcDvwYiyv+KS4TKEfeDTbqjDUszLuzrQ+
/+lvh2LvUMbioE43E8PYEbhxl8MW/fjj/qrXXThadK83pNWMhUEVQ2S+PEbym7BeHKO3uBAiZ/dN
BB4LpmmFEpIlA1zY9C47jpHCG4cuu2FUhuivUWkCbdCzZvGquRcl3hM2EbBPkaajPM75+Rfs4zo6
HXr20Gy3goffO7uEIB+NomSrUc4TSv1DIQzsWNWVPKCXOgOEOSTIJoOlV2GpPwL240L8h4Iktkq2
ccetnFCCvLuupcl6kkJVajOxB8CGWoZf0dhSaqXqNvS2rpcN7lcn2ccuJP66GbsqLh9AtiZ0nNxq
R7f+XIOVzW8S4XfoE7XF6UU+JEFQU/qQTBL6DY5jyVhh+qUroriFn5C9HSLCLSDxpPkR8lCd927c
5fxduMFxSosn/1t7XhFg0fltdKPuHDfwyjhA8Ge4fN4+apRuAddXf63O2aS3z/kBWGK0QCdgAIJZ
f2/9MIAm983SOvKvgTJFosvD2ZkKbrXaguBZpbtvziuqIrTthD5NQ9U3E+hEpW91Kc+J0gMwtplk
2EVQ9YbLsOGrDbAgOWBUiB873OQAyIako+N2XKWZOa5DpY7r6NPodKF2L1tI9ehptDEzxzS1YN1e
i1udUV4ruTptjpaGWM1UR8WMfdN8nrD/izaQWl7NqhD8YybCK4mIsva8X1dYalIUzs/U6b0ateAI
nAoG83vmQi9AWCq9oNhUvtwFyvSqHXXGTKwKY1LfNVFRN16MGauGpLQDUG3w6Pp1YhDt7/xkmWj+
MpKIbDBam8Kx39FbRzYGrCBecZdlGM0GJwYAcrV4l8GO8U9Qx6vUFJRMCtb+huNg5wVZd4xBCwGG
dgebjaaZkE9Tsq/ms7PlkeHtxoLlMTejO5UU9QzJ/zv4L1pRUKrHQQ2iO6ymAZOcMmWKiaZ0lDzV
ehsrF284dVChbxIgo9wmDh7M+68ZpLfVTZeDqJd570CzBLGO3Rv8l0wXzFTh3U5z7iQX66X+fZdi
VQq7oP1/I1X71H2h1g2C4J1sr7tEX8jS8ggR/4BOVTqc7g2gOS7kLrD1Zqgubx5s8pL6+6MFk/uQ
4qv4/HmMjBgGrccvriQ4H1eh0ZQSpZpx/5suPh1MzE4w9Jb0HvARPorkHNXhaIZv9o3ZXb3y+U5v
OSKdsktkDsd4hxy8GKwsAZ5P8phjayWfG7LWTnHKp2TAHk9KfPMpZ+TPX+5b+Kt3osyEPozu+bKx
2fzdfr046hMhYRHgAT5e+ZCQ7x5ejUPOi02mlbfjN8Hd1437PirpOYVJdHc47WLb6UgDXo4BbzSC
VTCa3z5xMaSJ+iDjEDtxVXIjaiQhil6zLcDI4NwgW/sTSZ4w6KGZvDsuNTlAgY9luBLbtiFUD7+l
g77vdm1gd9SW3B0bjxKA3gqiUKhF5WsYNbC0OusVjaK9gRVwhFyZbi5++T5bA5ahuUTE0uCow9e5
9faj5SB2LcG9JJJSB3dbmB5nm+1z+K6XspJqmfxmTqynHZoEZgA3pHee3o/6SPp60rYDzo8f9SB3
RDpnG32mOa5zTwolqhyf+6qVm9OHpaMIYI3qQfIlC3EkOwjqZFskSUWfq/tVSIU2kgWuM5drV+sF
gIOsK8rCUaG3W2c8UabGH/8o7bDDmpI7S4R3NrSCT5qhkUw8PS3f7fzhVlPpQdb3mOGE/0UITcsf
h+DsJCsd8seVB+FeeyIO4IkENeaegMJMhr+f6cdxpjeCs9i01mibYLdkD/iNc06sdXpzvIiy43TW
xIl5WatgrHgngC0cZ9kcWNEp4X5XpWRs8PQ3SuAYjAitLaAMsY5DOA4Aw64TXN/0um6J01FaXpHf
74to5a+FDO5R3Pr7junU6joFzRKsvH68wSxtdr/Og3xerSjTErdRmw9aXD/HHM5kJ4p9lrww6XhD
kywB9U+cA4uVDBCP+k+BPIOPBJEhZbPLLXmMQUK1vcrLUJKkJpWodV2JhppLxiPfeKMpOyFNx7F/
DIdZSERsATMhDtrmtbiiXeiWnlZyxSZsR2b0b5RcYl8eIvbeOvP60Tcl/zzpFtbUFjVRLq25gUCD
Nl7vhU++4ebs034/lB0OWtVS9jD12Ncu0gpMSHilWfu58rBoiKHgJ0Ixm1TfjNK7hjZ2PygIRiwU
p/dVE5qC8ygso0TNhgwyEovqXstzL8OUvpQCIWCyr0G2XYD3ZjX/76dK9brCNJkZdX+24jLKC30t
9cpO47Rk6lHXV0PyMfqD3swDBRxXrwfFmSr3F7UAUF+o76MLTOUznaWwgavV8INGA2m9rb6uSTqU
iJwT1d0GqF+LP4qJB815j9FnZmjF9TBinBYd1AS5i5x8ntpHVuwPMMUlScrE41xX9jDOAhJh0Ki/
KJevdOSPew4r3ty5cRcd8034ByQXAnMRWi1M+4i0PrNnJ4DRcuRj79yZK+EuzAtYubGdDWMFES89
aSqDiGhiCFz1Cz3zZK5Zx+zNYRlsV9xEuhlvQe1fL66d6LObG717POj+ng2b2h/1dHEnZTANnBZY
iE+kAZFJPfX3yrqzjv6OtOV3gO7U8Mc6qezF0hVaQ6l88P/dXMDoOByWfhtsHF0LoCamA4yRA7df
QYY//xXheuUSYMn+Z/zKYdtJgEaZqKNc6xH/tmJivlO9lf3w2aNl1MaGpKDN9WLwZbdiaXdk+VnU
AdetGlgBZQ0HnByCoNoqNhgQ0zha2mxRfF/Dxllgj/eVjDn/owDZFXUHRgIH2SerMRd51RaqdoN+
1+TZZpiRnx6bFVvPQTvRTh5vkaKTGb6lCNDiHOMJmracl4t3gnKv/Vay8IYg5EhGpXlvATCr4FEl
OjM85HDzd3wcXTZQXxUnmNx2YJHbqwKSWyQIabPVy5rMG8RGPFV4JPdHgRZEaNA5p8+/FWfXG0dL
7EZbpYgaukxqQ/4xcwIxgufXt/gd5kNRzaD0fIY0dzVWe50GnJnHx37ZsYTxJNdQPlGE5PpeSN3y
dtTPtdjHgLVFPxHuBLPEKsdlMLpbFqZqP3eFjf6tMp6zX1paVUxkkz3SOpVBGUBdnsq+7YNpxEb1
B19JODaKCAwfwOrl0O/wYjGNi+fvdmg3eA11dImy/aU3HGuCGx/4FwBsQErp+Kv43pf5QH7Dz8nb
4ffn5wRm/lQfJpqy+MPKmnPK5MebFIS3jLwSus8V8hVyHdRqmwalG0da5eDi9zQ9hV9N1spVcO8w
cE/glK4YkLXJQgmhrCrIkxciNMmFbY+P71jEkUCZUYHstGF0CoLgyOTrB1WptKXQAOTaqw/jWIz+
gTwijfhtjCF0TG2P6agelLYGBpykwVpt8uCM3HptBg6DSPBPQMTMRIGVfqh3Zvh8OGGa0jsZd1tk
dqIWPYH6SfYW3O+vuVzcEIc4gklPDSjTwVWf6oPXDNaXyPqGWXLtcrod3/3PCg5EaXMzGccb3mly
pUiKZMvCJ5VKP10phQe+l8zMhWK2cvBWtZJ6pEhh8awUCiB7gNLNRKidlYwPM0DP7qTKdAsPyJAk
krbLo3NmI60tHbweJEEWV3CAsVTkO9vCmEVHvp1GI9Ak92WYHlH9LZScXFgJJx1CwgeS3dbIVObr
/1y6RvZKEA12P4LBBq2yCNZ2pkRmjMgXrgW3abYVZvJS4r6nlKPD5xPjv565WC2j09wZ7uRDgyNR
yxuld10emncoH6outZX0/k3voKGM8gFgDuS/aH+o2pX/Hr8K9G8JrtDpAaL8nJ7KEYyJz9kTQpVR
Q8zqNgtLAUPH54DVWNnyCIC7oPXUBBKXK9dJfScuJN0QV6xsypF4Iw3Px41jMARUViXvjY+0Eayx
9LO6xEwBK+E2zz1+xR+yMi6s0FhdQFOZTxxoRO8dr9IHqW50Kaap6dIWuYJtstd8T2IhXmU6tOTD
OcOu+JdThqmEjJ6t7EQEboKC6uONWvAjUMdClVRXCBXKZWngqOoqYq/y1ycmVEjwxBdOm38DgrK0
8kKAatAIoFPem99z1rPXGRsjlONGa86uGcSHPyKtutwvsJv39bR549mMq7a+sFdFEQT6Wl16ZZpp
/GsLljp+ZkAp6onX2qQabIcu76gKbM0p3gu7v5LNEJ1phzu7zzZ4ZMQ4zWSCUtLZj8HJxiCFb4SP
xGB5l70lG5qKKBnWJlzkbwNlHHRMqwR+c02oQVChmWmU4vsrVoJ4bCICcIgNfC+uryoMRely4xPS
YyNpnQwS7ttjTO/NAoecouAla1F98hqGZjY9IR1xhC413NQZY6SCJlEzo7olVfTLaTRi/mnMHLOj
yLm9Hl93NwMArk8q95sdQ92YkoA7RU627S7VIBxQeA07wQcynGoNwf+GIhdUHf8krof57j5MtO2H
TV352vEH8Z2UiIq0tafd4c3NqkIK/sJXFg1C9bv2n2L8/iNa0hbzHI/001j6v4AZBnluZzv9qvKp
IOSQKB3pK2nyxOU7YLK3tXHUsllx5Bc5hkaj1D7rWHRtng0WM8ccqitaE6oLXO9x9+F1YVcOKTKI
vGg5Al3rXqffwUpff804d9JRZciUJxTkgvNoP0CPnM3KV2WX007/oJfVbH5vG+KDcQ2AWN2ldYCy
fpWvlmdJBY8s4LSBJ8MCAZ2mCUWrNWcuRVzIs5ZQXHh3xzUvTA6fRyy0/RIRq2kR4bm0qr5rXDTb
ObLoZ0YMterUE6Uex+vVMJisCP5QrYmkcndmddOkcESRtyDjZx88VKbW2L+zW/AtPuOkozIBn9hF
wKqw/C2QD1BFFWz2BAAWc2BeHfigVQynzkBgxbrmAetum9rOttRnidvikdsf3voYSUMPjp8+NSdQ
P8DPylb2GW6a0b9xrgyaq3u176G8K6qTVFjoXSY7RLL9/9uHC5AurJBFVtsQxVxbQukiEUeb/azp
fwpGo8TNdNLbU/MpPCgQuc+01serw1aGg+zMUjCHAcSi7TgweECsfhElSm8XTbOykP42BWSDUqUI
uzdg6/Bpu7679vKdr4dQtWe4iBVLK7gvBXlHzp6wW4axWe0XLXwr2VTTHaR9Jl8wWnHuOk8tu8ba
x8B92NK9LZigaMKyjtD+GkYzTIYRv8xS1jRE2sBsuFYW3BokzJ25gC50WL6XgZLnOnslyR/OENz7
AGI3cXR2njrMW0cenBvBy5AoM3aQob7xdSbYlklNoB4hPqLf7vg223R9dTfEzMJkQM3DSYuhWjQC
otyyCUC0p9DZh6B6SwYE9bBO83V6wnGGhsCPDclliAK3/ibGKlGt2yZ3A9NN+G1m2b23nczt9XBE
aPz69eAeI3h2iyLs0Dsr0A5Z7Hz0/gvFWPWG8cJOJ3CXYBv/R2kih8UHJ4H5XoI+au+kDThdBAjW
3u/ppjQLVFDl0VhWcjbK3HeqxsBMX6GY4tbzVAfm6s23FpHMmBzVYZZe8jY2JgPmyzghmcRoO4wO
FH/e11/J8M1G25q3u2H9Bp2pTo2Kg6AI9q4n7RzahZ+IBX26HwW2avXk4ibjPIc6UbF9U9fshPEh
K4bTpg8GzmPpLeya/YrUwAMtiYO38HxE0881bZyRGX23uSHwW/UAqtx88oUypTqGooLknfS29jKl
2Kmz3PtJSSJa15GmweybiLmSpVp7rlpnT1VeMfuSCarxPOk5C0w2ylBbrXTUa0kWrqhAyMLs/N4h
1EUx/cQUxTRmeoztbet27hYn4EpfYs3hDJ7R5ZCsra+YtV0ksjLzWIXVIZH1n/9p83wYyXRv8qPc
4xUUIr5zZnJsYzWges/9suOfzJhm6nVyH3N/F9s42cBjjMAPHJWIhCHjB14LCF8cGH2eNFqd+glG
9kBTuljMAPltBuVY1kEtY3Ccpm85N+265srXIvZluMSUDHMtbfoUb673iVvn7kHxLYV335QUvMKO
aDaSfX4ky3jyURzJYmCHLJprhlXTGnsBV682J+wzihxrWEnspcjHr1dHNgT/XMciS1z4ngWZti5I
jF+ZNmt5F/O0D+UXY1D6aDNoe1Tnsek+LzxYDEHvGj9edTt9NCIklVqqLRrQKlB3NWQD1h2eBSqM
9BCwBM1Qp1xkpgnu5QWdl9lEB5Ej4XNXCyhoRBx+O/QcPmPBoN1h41ke4CY5LiR+sIHjvbVpQk02
M0FpT46AmbXT5Ewfe/XGWNGsaM0+8aEQwQdmgTYCTxg/cci6fbfQiS2vmP6ztIxDd1oYCPlIXAvC
Z4TSPadyGTJlTjLdzjeyuD9M9UI1XOgICooHtzzi2C+WRrozssIHY3mYt/SE4s7qsUV5cLggg/D7
YOzCfQd4SAOakCc+n7FRJnjpJIIlgvv3LIrS6YKXhZClTvcHY2K14cKLClH6/qoBcmEKdHbpJBbA
lVPYIVkNmXHFyaJsdEyahT0Gyd5T8vzObfqZw1CFn7nyrtH9WXZhXvFHUq5RgpXHfgEP2iS0sqA9
ye/EjdVSiOT5bB7zGT4JyGMLeFFhXpKDRiLMCR90sOJ2eX2d55c8sN8b2UJWzWj7uJm81LBGrTXc
yJaEvDmcDyNFl1LqC9nzRvRTdCDqVrFhDZXve5CemwnCHgwBqMVFcAUkAdoPKfszNpYwI8c8LQ70
Xkrj0vO55b5ZYdHf5ZQvSWpkifR3O0bXKSCh6TWP6nhgeVA4LRIeMzdNNrrfe7pfekSOEXxiCL05
O8ubB08fnrZNiYHLsE54WQ/TW6ptQTCkLVMu7WWrMO/F+yypV2NFfDChIPKoc4+mrdupTXT1HJew
IX9g6AbqOEGR4W+djqD7xDJZ1+CtW9u/RvJlVfwBOtyG+cxIW6sqr5OWgck2DrB4ZfzXqyWRLuZv
W/fMlmTspkfi0+Z3vtqLJt0UAvUH3scR/fT2taEOB/ySZhvhwTTaxcjwFKCi04iu759aL61Ujpz8
FQJMlJPgfIsbzE/Nv6ep8m4GMeVbxMwpqClnQl06R6qJ4wjSt2guYeEL9cU4TkNKeXulBwbrtYtO
QuaB4kpnFSEm2wBc2X3TF0U5RbmlySRanVpHoZosx/6d5zDg6VjhF9xWZALISmtgLSsXFsbvwnPq
cLCBIS16WagGsNMDKzFNTBrSuLZBjz2bC97+zYv2f7k1jY6Aqg+s3Zkb9DwXKy/q+ovNf046/edN
xU7uNcNGe/jwmvnZ7yEaqsE3uJNORvpKRM85c2/tm5Cq8ewGi110dyk9pPtlIUlSY343fkdq1nfm
2MJZLNgCONNNaro3sd6fS+wC13ZzIgynvTqWDyvhRaItfEYMskL0Ae/IB7gBhgYYVNHhVomhNQP1
Bvh8w/f0EgX7kj4jejua+o1/GaMljyQPVCd3yOEQknRBs52Iwkv/ZZpqoXmnLJyT5rtdSKI2ExS5
zqyCqXujk27bZ7VCZZ9WL1AA5KITX917cRLCzdvW+M8zJA67z7s2dzioGiXjHZBF6IomqPIuFpu+
2LvxbMEdkQj9lJtiaYBtrbLNPA8guPm1NmMXPerCLXtWw7VQMNz8pY92Pm4xcu8h9u3OpUa47vGR
cXJFn9y1gmoC29ZBHS1dKQSzNS0aEYPK0b4ZalF3pGc/oKzlHuzFrZmbXgQOL//U2QTzkzgdNzJx
k5WGR+mJpLuCL1RYWLMJQwIpYQxH5+Bnz8nMkFYyH8//9PPmB9ToKcAp49E+QCRVz0fkZkDbtS1q
s3DDq61E/223D1erKzKPw7cB+tjmAF1yO5eqt8PM5yrefmBuoSqBJExhw4Isgy8uZ9ne3lRyQpZ4
9IP2zYJlITQMQa0STEvLAXP2z8OaUrmulOVTheCt6bA8REnY0MeRuyjegucPzA/3PbM+dTbB70Pi
RCFeS7hp+od7MN2QGJpCOTr2IXwexESp/Y9hEvHw/KOdbQ7YOktABTtz+4i6n/g06s++kzhl5wGu
Dn7GJFka3alF48iJny19qhzuYl5jsW4kd19VS8aIvwjFnewFJanxqAcl5zGy25wzanM/hXWyICCt
F0+pK0qiK8QWMU5z5+9dp4DBung9fHrSPkpL0fqrIktgGY7CiYbHd6nGyKkUGu9B/Yg8biZ2N4pM
YjUWCAdUSNnxs4iDQ9U/NrJohgdgopUetmcRT0scvr9cYEr4k64L+W3PkWEBNeyLF+/XhJaQmC4V
BfveVfJ1vFg3hKynJzqOl2mWE0Tm55ZIbgLIiq0D83L38N06astsXu/JOUiBT4+mnpzF4mDm4Rif
86SQe/pq3kXuazEEofbxSyritfL8HYjw5kQquI9uBv9reR84c3MB/UJJP7K2GNSIAniKqR/6p5c/
GRIMhi6JUDXGa5YwXdw1cESGMhBDipDv7heEjyOU09a2JqX8Mx1TeG6rFMfeceAD03lxL5PY+r2v
uqsQaP7DnIflZS02esLoBNycSF4SA7Cg32Ecz9uJqKyNdfN5aRzcybq8YzfdgduN59PEU4ojoYMx
i96NnnQYWzh7uF7iPgQzYacV1cz8sbxaBgncqpaHtg4KBDaCSvTqs4NbmTLUATOydtPV570oewAw
ZD5Hu1YU81x7eLh/axzGY9szm3hhyogd1BKXZljo/RZ/d5953/RWpeJ+1RhoMqXrd9vtNC1nPtge
JxTdOxkf/GHlUfdDhhv3eRe70fizlGnnsR6Vu1oIiFB7/MrL7q6P9jp7TKVoMp4W7bt322LP5Dqn
C6KpL9y47NXL9LDWMQxDLzyFbV3w/1TjayvEglB0ifDXgYba/rBmVH729Do3NY05RzUhPSJZEmiU
h5RXSabGZ2hpDsbbNv/4SaHzK8/i3IfK8xdBGO43mhkHhGR6UVnLjA2MWFT9HiGUAKtqfLPnENAH
j+ASJZ77vF4KzNxCRcMgDhlqAQMENIOdBKzg2H8gMSt9eV2zJPAIKhtaVMgMEXBkHUvGhZR52kLj
syA5uHaJ76CYXnpfk5wxKTYHujf07ynvoMmLU+uspHDu3cssf+aplBXMNWfnnMXw1/l/ckmz+h7n
YHbgm047FozBwvpndsFS4zTOShBFL18i0RjBw3+3XrLfJUegMFrAMSP+bOUraMpcXF/4UPGNlb8q
jZ4/QB00/jNDZ9xGF4ZpZTySJBSshJMa2rjAIUYj3DGrriA3livOKXKEFsSDTxE+f8zg6qX2jowJ
JZ6Cz/i2Bl9bKsnl98190ZuV3tjVrMu8drgQqwrxdkhJkIZC/CDa+USlvU/wHrVTCipHQnv8WKlk
NLY54IbLFuVR7BW23qN+zzasuQdZhS8xNt4dvQmSRDbrjDUgwkj4tRSzc95yK8bmKjkeSWF5ht2u
v4y9imgDeSxiEP991PNrYJ6XOc2KbSR6W9/AdlyD1X4/2PXYZz9ATzs5xts5Nu3W9KI1dNMXcUgl
5PixsWe0YtlDN5Ym+zWaEMG5ZbaHcTKddMN1itOPgnMF6yyzj8LQtmzjLFi3LeWKCsjkoYPLjqO6
TqukayjlzMajkd9EcVbKQiaeB0JCh/BvK2fiYq6khLOUBEMxnKzd5phhXI70KjYv6c4BvOPwbP8Q
eeulX8I0iAL4cVWclQGPTtg16r05BkXPi9JC/8tLQyD2dnvkQQmcH/uK2a7PTpo9qS6w17Rb5WwO
C+zlQf7oAtMA5eY26i3nMmjpFZacuIfEcDB+0UUdU7mrtrCzqsl7Uww1RNdkywP0hjbLK4sITjhi
yeHSyEOhCYGFabs9+VeMaXOcwPZQnpcoi+YpY5FWcKNT5KK27ItZGxi5RdYqEXrtgNMvQGLL/Vgw
Ik0BCBJSUfLEfOGH7cmtEMFE+3ZNEg63uSQRBoft87O0I3hDRAgIPHJEh5Pi9TOmChSBiBbav33m
CXWCJ9/dbbVjZxWphvaXc+MuVoAVCY5h4cmQv9P+LbHbciQ/3OljrZsoxZ9+MgiRganSnBt/7/mg
jQ9Qs9RKQmNfAxKHEL05UHHRPlAuGBJqEn+kxrTEUBfLZRbR4GcqIv81HzGlq6XMT+whClBOPIWq
bOoHX8NAUnXWGdgQn0Ju3Zh26TXOf2r8M0kDj21yiefLliJdtH2+IUnrGVByG70CV31zC0nY1VWi
fkTK+cyjIeTTHaoIiAo8zym3y1r97Y0iAu+rBcJmrX5uQ6o+pwXQEreQkJiHUZECryWeLWI3biVJ
DDq2WsZP6MVM77KVx2790WPQsBbfJjdraAZDJl5H7fswkJWZvClIEsQbHg1BeeGEbE8Hc5bQ3+uj
c7vfVYj89NgeDIH5TUnHS5M0/dHBDnlkvVRYljWXvdXatk9ta5ucHICOdiu+ODqMV4Gq6P8zvQ9g
T5Rsd/aJhv7UlztoiX724nt9DwnFdKnJAYUpVUgc/1TGOOKzmD9qqaTZYzulhuBQ6V12i0AekVHT
U/GlqMwrtKuDXpo3IXmHHOWtVNicc6n4szgY0QJiSok6YSugbp/EB5fJu11I49akWuTJJ8CRRv+c
h2D9UoaCM+vsDUmbC2vtyvaOysS6ixmsX7NCX4Q4wojL+29hfJrkPqdlScRcAC20kUi78e83hiqp
9NxZYh/rDm70D2Wy+3mMCM06BI9sUKkzKaJLQ53itOxgtGiLCD1bEysReZzrC4MPqc5OUHO0l3iV
feGeJg6At43z0oOb09VU2LWccbP7A9/JMCJ6gPcuI+ZBl0fpEIceJ6nOAmP528lRzPFdUoRsextT
s2WHaKs/wfJ9N43GjkT70TM8jrxG6/AJyVu159wsBJymQ4o7QvH5WANyqZgEMoL3XENx/u0wMpMq
iQyh11C+f2Wm/6uVCBaPeUYjWjOl66y0nmdSY86fLrrRNk9rhKMkQfpFpXpGGABgnv5YG0bP2euF
3cayL1qG2oPrHBH040kGssJPe3SK2xJgTODFTeAzKyfmEwjah1AugturRt3aOVtySIifmmPzJzgY
zaNouGjMtpTyc8SfkDBCBtePrsJDGRKcjGO29Z2trJKoT/kCzcG7P8jp4p20nJYd02rJB7lweQ7A
IZjY8hI2wKxJmwJk5CAilsEfBlmOmqGkCkMd/freO6XNIYlnbOG2tN2Pj4fYU3XBzb5uD0HuhZEB
ZV9BY5QmvGqgpb/tmyFSBckFk1uT/Evx394kVKwLg+yBl2Y+9JsZDzelqKsNmViqajda5HlyTPil
mmhB+Gg17/ENEZSg6YCx5+zoe7y/dd0B9TZ1Sfclw2lExmwkMN1BSERSz4VrVr0hRtfL2XYDCQ0o
B3zWZwBBD+NHQEACZBLGlCySl0NeQC6gn8ci+gEfrl67oKE6gzjbo9ijqVZ2sidFELHcvA0NszyR
DNRsOnR+9ZXvmA+8E9Qas/iMGXMH3aktvPoP+SjDHt9unAx4cZrJtGOLxcJNavDVBnD1f+R8dg35
V6WYSHRQsqWlTtP4Q7pmzasNjJlA29lK2IussvLti/G65w8yyxEhOvE8dDQQVSmlkQGlOHQGW4Hr
x0ejGr2/ePROJhTzi2aFGa0C+Ew6eQoJTujY2tXZyvP3fVBxO+kXIwF7gSIoiq7kC5pCgeHfNijX
L5kvu8EVE5lWhs9xrENYUkAKoSZ7ZivkagR/JVyUjlhPFuc5Zp5QqvnYYMEYD1Lgrb11MFm4+HAA
fsKHPV131veMybNLPQW8SXXWwkByq73YQSxE0NLmXcmcFDAxyHKEe8bLEoxeevoeYalhasqNfzxO
oVBvzrLQRdV+IAx+ECQLUdvLH/QvDy7lBnRA86kKpLis7/QfCmW3E62O1vuQz/Txj+Wjz7S+5SsV
JX471NCUCmNEWlIyR247dvnx7LLqIHNc8e+L5mpR7h0Cy8lsBRRSOszbpsIHQWyAyTBo3GirmMXN
rJJZLLdfKHE6Vd+gj060Uk2QoE2uFVv0PbXk7JiG23DDoBG5Sr/awNO2wP7nwlgtgxel17PkkAP5
jOeKzcs+DiwSSAXf4fNqchfg5q8J+YPq8Nbkdp4UHASlN+FyrwTmsdMwuF/YVJF8gcQQX3aJKxte
i7OMmNJycyXjZDsPiw9GYsxVb0ahJf/QSObNoJsFhV5LCtq7sfXhjJIFCLFpuo6LQ4EsYl7Pyx2V
i2QaLnV1QQHohYrIA8PpAkwN1HbMZBLoY7UT/zodoreENS/SzeQMlCpVEdXbslBvFG6nqE9BFMmL
TADXX8p6eZbeRlnYgUe0PrKHT1BvjQfVWJIzQ3B3JKHZBwfv6m8NJs84msrnxtWR8yxdkKA9I+x5
3rjakNVsjAzAHkrnAVUd6kEdefXu6nTYSyDKdcchTi11XpsJFEaR3nUmerUE6HLeDll8NelTByjL
J1YXgyXm14mqQ7ZN0fUHQRJLSC6HtRDZ8ai5QjwA23Ik0Q977Xv23L6SkiF7pg5SDem8oRp3q2Rq
TXoxAU6J07p/+Mm92/vNOgsE6wVAQOadg4YN3xGu8ZX4J2ifF9owUYJEU8jURP4gqcLFiPL44dYZ
xkv7mXshyqBTseX4NhCu+kqvu13qXHWheZbCaK2a4ClNuPYOyspvD/MRwHDX0yOB7onzLOFLR3bt
IZPfMIYQm+9okRQJQXk3rzRajzYPs8hYP3ZxLpY7fl0ZEtVDHvycKvIgKcuSO+CLPWkzwuCee2UV
HeEnB1SSWNfaPmdWn0drGd8vd+WjdfQQa8puBxGcDxS+KxmZrlLX7e6+dzr+7IcrN82LlEuTZ3B+
FvGvv5SMLyeUyaI1rF8v3bBGe8ko/oNXlRt3wkNnJigmgAET84UnAt63DDFaisG7YWd/TlYc4qQv
3nDUPeElAlDIPT2KBaUZQIl0Vfn1vqvdJhNrGjg2r3LImn0Ioifw0bExHxqxALX/7racwO3H0jGJ
XbP16Jo9Yg+MlB47UjGY8QZJ2fl/JCjA91UyIPsdQ309R8l7UAzUnrRunrFBbcRNnTQzCGMZ5ug4
PeMsHpXa11wxsSrRLmOnP1AA89ovSYjJ3TjzY901/lHOrQ6yKhUH81CP1MMmJ6MvYDPgE71SiXdU
EO/4Nx9a5/hY7I7tTBTJf/3wMIKf1ZTcUU6qUM/Ddf7Rb0kUdnJeEjIP9M0UakHuVv0j9kvbKaCE
mQxf1XNQX5OernBGeHEZan3vEZ9jetLZzDEixnZbeEiib5WP6mq0WRzxdRgh6zUC/6uexaaiBrGV
Ip041jk0lXWi8Ayj6/4k0GUeUdKt+SkjM2BZEvQBEttqdFQKpW0piU40JYICwmqTEwf5UIHF8+VM
88I4KKVyG0XxaL/ZCMD+UYks9tOItZbGr7rpySUyRkU0ye+uW3hKuy9+XCY7a7zZPt0b+8A8KxBq
HbvURtsdZEWrCrNC4ihYMc1wOPMJFB6axZiqkzqesjhQQVqsM2TpjwtC59DF31CvaJ1pUcFoI5Il
P4qdIfgb+doFyzay5mkvo/WCTiUMSEZ9kRygqQ+qU3IK8NR3Ed7ViERoMiDVcxvWDKjmT8/SkiTq
F3s2g0MhMLOhro115zUzU0Nv2PRGSxgrdLshmOar99onU9Vw5AriAZwJCapiWWWYnazaM3lUXvI9
cLF+rDkZue21LnHzSaTvcw+bF4OXjq+9aH8uTtlnAkKyRF3pjYk5brfCPHQlmlaz0tX8LTvDWyWI
Yp8OcbD0n5gsNlU1E1GKpx3FaEy1Rh1Q3i7g7gjEFk4ttBAbeGHpH8/3kjWX+TxGNV2HZ2W/EWJE
T5W5/UZsOMIyjvMJl07QoQ1lihsIERCR80H8LmAqpLZAQNbhZxiUSUdOXZtZFFejpFKqc/BSr1ni
VWemTkj2M2PGJJCYKqzj/0LexQwLeLTbKKzl0iHwR9HgV1KaepWCj3Ns8uBA990E9mgUzIo7EiFP
mI/fws2L0DxxixIyygLTCFPprxrv5Pt4R70a8yL/mxfhCyoz+PfGCEgscCG9Gq6XULRKBGdxEm/o
UreJ5fpiyhovi5qdj5eAkPUG+HZTdvuBohBa1a6UP4jbdHzdWgs3a8BM3ox/ZAvZR7qiRTfckWFc
YB5KvPiFnVMgViAtIRwDQVQ5bMp7Naabj+1nUNnG0e8jPY0SDBu2fth/H6sYsbP8nXB4vCQWQOnq
6Gdqe3eP1ncIuYGFzKDFrx91VQSHYr1MCFu7HLWxMvNXGRRtVoqBLJz7LBL/S07iPpcFAPbjGAKx
4UFf6xESzCXiLX1mFJoWpTTYEqVHX/j3TMU/+0nnC8DaygvYwEkkq6USta4vxxRmr3UJBBjIihXd
VOXrE9+84hyVyhNhKD+s3CldeVII+a5rjKPERJ6qorlfQDRDtk/QkrInXNYMUzo6J3jRYPLsmg1S
4mQBkQVuH+fU7IYJ5DyDa3bwR2xYDdbgLh7qV6nAZceAMGyBANV/SjfLsz01rBIrdmuJTj9N6HkR
+myeFl0odPODhodNWTs7ElZ6an+wgzqSlDzm/fAkyWGU8QgLmRlz7s+3Dng3z6GBxmKA53wBTfNd
4TvTs9YXqdu+L1Zp0RhGYf7IW7EIxc8goPGFP15CcTGaIdKEIpDx+M3avCrk/dztGroLWXxw0hVP
pLQYFnbyN3CaL0TOpyYUTyUji0srJV/497FxIfl/kx9zy+KQ+l0sZ06heZiwmD4vMnCAmgtOGHN6
Ac+M8fWOIJ7YSDTv4hB4WbTbfiMTbZI0HyaFOpLnjIxvA6abi+dNo415iBN5WkIbaHjhRTGMmWAC
Ac3f8QvxwZN6oj6MA4CHgsZ8lz87gtKh4GpaBqxcZwj+nbuIyCemuCJHYqehEXnHMkJa3hXJqpYq
YIUdW1psBlIFaP85q17/HWVjA26wJyEX5ceSd5rW/iPZWScFyHsotbNlBkpJhLJBrn3XJ3AHlvn6
T6f68Nze2F3U5xZeK2EVkQu4vZh74mrfJ9vrb0WkAw54le9OWP4TNZ8PMEMefGMg3VPF+wxaKxku
Y7mcQ5PuQmfIvN642diHDk6BNveQRDQX9Yq8NMl5Y1fFXP0500SPoa2mtdifsr0ZTRm82cCpdUYr
Q/58wUnvwuSqgCCh27JZNYltwCsinCSO6K0vZh3ez0WB09syutY3H44uOKyHZMbuk0Jr89HM60sW
CZY6lym3u0Cp/vzZnHZvaZkrYsydSQ8fMCWPUaYNxGHunRvwFb8gWYsKfM4B9r6C3tqvRwYp6QFj
cHNSVm4B+Rh8IvTxYutuB3MP+lIr8nbIEaYJ5QWaNQZS2J6rRVdQ4Gh+B4C0BE6i2lsePO947TUT
VCW48mVUnK7IWw0daXyQ5CIES1Y1WLbj479qWxot3co3lN9hitFhvnHddksVTsSidh4N1ma0As8v
0IE4brzIU27PwwuvP2NzxGCEdlYlJ2nsU0cMuPe3lISwqRQTqHrRqYnbW2iP2lqfxXUgIcebhzuf
djaz4zHhC1wDWCiJgWzK58kwQMJZy96JMn1uZ9iNY6zfTa2fYavRV4Fw92TBejxZVo5kDgZlFfe/
AKfChxQi8VwOte7u2aAps9jSdvUWbYM6H7mF8yOTnNK4VKXPlsM0KtFzirCx0vSdgJs8pK1DGYOy
Xa76KDUVykV1OXuYcyHCr4qJ69HMpsdxV+zz/9Qk+qwMnLqrzpOTvImYsg+4OZo4HM+2hcgFAoxr
OWGXytSV0UiVo9SpqjFEjRIkjiARmFC3U7QCo1wRAYISp4IS3RMCJBc013Qu9/pYLdyqJ/Utolt4
b1/MmYzwHs6PzNMF3lGY+AY6HcEEXUqBb62TAxAb/5tO7iFLjGpgG5KPDw/8juYZlJUrTjqwjQPC
VJbduCHi7xWcPQu01c6GbM/T/pl+Js1JWkUbYMyv6HSUb2SQ9ecaIyse7u5sEJoFWJEdi3GD5Z/q
QrfmLqNVg8raJU68B6nvvGrRFvY5A6gN9v6OepXrJh47xlX3RVs8zncoTjFKaz4dUFwPsN4ZripU
kLpD4NPZQfwLwzHS/K42TdnHwbzL7Jqpkn9t5p1ceYEf1SJlGhOUVr2Lejy5jlLIPZDrvhmCpNb/
YkY+SjtX3lKxS6294mFMu9mSFOeL32Lcy1XBZleGzuLSgxKoNwYaN0kiS1aXhcPqKGhUWULcLgWU
3DkHPkCwR6NG8XfPeP9iYSwc5V0Dkfvttim/K2NJ3qdU2+POAHInCLW75QjLR3UaMwug7UqhzgvT
fMSQDV1zWATWFDsOk6aweSY4jeuxwevqMwTJR6pmNb5gc0amTNLDVRQ0/UAf14z3sEVa3d40fPt+
X2AIEiesRW+0KPLU6C1pYZxD9IjmTSzUW7Vtagl7l6ju8OPlwib/38zbiYrXZGBthpslglnYlFji
CyS3XDVRniOO0DJt4LPphwjgELz8nyOnS+oSvWQyic5SdqCF19dxqvNbwNI6CXP5ytd7kxwByQu4
xJjD+T/JC8cb3DUvKHBJP7DueZjnbnlVZiybU7JjXIVh3EqBDNF33Ooq6xX/pAWisI0UVVb1vhMA
6RNqpeCYau6GurAXJuy6Wsds1XSNKpdEX8/+dzsU7V43YX/R7KVQf32cuzotiq0A2CR/Xju/6RdA
kO8jgHH3qYIemMHxKt4x8XFFaeQR1buPIir0uDQnbn63y0oLyP4nz0WPLCISh1S6fCq5xNmQaYw0
UDl8oMmX/PMr9FnM/GEr9Lf6laFRLIZF7V9v1iyCBdemqjFHO0XWHz/9c5MH4PB5KeM7lFVRmGLC
/iXTVsyF7U8UiAl/95dOlkMFRsPa8bznBd6yQHw3eZsy/jKM3dTtaCwwV6dQY3xLeAO0jUJ2dc0N
grXl67EO3myb1/nkBwq92azy1neIZgOJJe1exW5ld1cKiDBZzyl7vKFr1STnFJmY5UER8GC37LRj
LHDB9kWl/Z6DY49RsMDKKQwglHg1QnarlvNumGSCxadMAz+vB40I3g6s2vFZKmzaUzon8G86BOfZ
KWE2NyFsSnhALVHG7KSw4BdPZdiv5+j8CdVdLgSmTbyikWnFwbCVmB6mTHHyysBrXijxmocXyQOp
muF6msBJnWgf26KEUPPReTQSFRwty9+qKNISPueZrvgYIxGu1Q3UW9OggZQR1IBFj+56XI9kyFzk
ypi1y8igVfB9tZmAcKusIKkMHKDPUa+rDPQ4XGR+/VxhV7/yiA5U3T2yhRGez3eEXmYuQ1SkhFuT
vW9AtX62mc4l5YB4uwjcFdB0U/dkudju1q+TMxqcs2dNvD1U+YwxF+vlJCyBmgQMLuNtLhcNcZhB
qq9cRmYxCG4X0BKEhTcY7UfwanYFOXyUnUQ/QOxFaDOeZ3KQzaKLRk4xfhMsBAz8rIqUcCq5K4kB
9v+bgvv4POMdtgJ0qpLbvTSG3og4wlRtlGOKJq9h1bciQ6F0Vkok5qDOA9EY22XQBypqMSc5rlq5
h4re9BVqEopuNG/jWE6ZelMMy2gTV2eEDg3lP9WlYQc6872EZBWPcyZ2Bh1QvDIhaWP3GH960R9u
aJ/8Sqz+rD1aaJk699d5gCpfxphBvL7B3IBjengvaWfVAH74eXKPyRex1ImU0/5UqrL08LHDYUy2
cezf1FExYc6HKIeMYn/1/WL5UyStvmbgnWCmmIQGt8cJNOq/Nb9sSB3ZVAoR/si3a6BdcsvuoECB
TCzhoe12LrseEt3x/yPy2S1S+PxNKPd0W81yryxQdxnJWe6T0B5MVUmSxqPAc2WXvw53Hu6A/ZUm
+hpaJIlSMD+ZoFOKhvljHW0rvyk84SdkM84T8Ld+zym6R8l8tb4dnLXauBWruYL0DKVNxpXibQo4
yZcl136sWT/yQB7Nmw8ZdXUzBLNtoyiyufqLz/9KMHxn/QEF7TpwAtZPbyAUJLc9XIcS2Krn/6Hn
di99Zx2sQrOsq3izXT+i2aca+4qcqSILfWZwdChpEHJDPJmC6dqVbUWN83MhmnnFVEPgBvyh9ZPu
U3Zhi7jEgTL0unxDV+sDOTJ2R+okUNkBkz8gywsgoJIqBF8A2uGGiyBQpt8KFpeaxaz8QB6ljH+8
c52unOg+dXjV82LUe6Kb4KhXy/KMwYzK10Tc8gdA8TI+FSeO9B3M367doaP+U2ZaoGHHdlLBo+ys
EU5yvl/SW5Zmy4rKvYk/uEymKwO1lVtyZCN/ShCTv9UAFZXEgXTs9qg45FSZOje8BeFyh1OlQzpE
ab5nSLWZ7+CMh/Zc18MPQc8XeEjeV7Y8BqDAgqIC/HJeewzCkXGTlDu5UVLkds6glaGNBV/wmQoy
1x8H8PHk14xSZNmSY+PQwsGPTbI9Gu7zaT8wUXGlWVu6nAkTO5wt5LyDaCKq4N0w5g91040O7VvU
k6PefC8V12RhXm8ozkKWihtOxlX4idufjZ1yDhNXe6YhAHKPKdR9WIINALLvqOU7YyG+DJ+scTdA
xTOOi3Ok6d+tpmQ51WJkyD1qDv/PBM1a0KkmY8ppGVKvTiRvYr89K7lloH0PkAC1sZ88XiuNOAEP
5c3iKIgr5d5Lruduf9hvHfnqbaP7RKN6MxFVgEB5eNwb9G/W0SJSYFt3CRZuskViwbom7YJX/VgZ
sB1lAA6YEu8fuStQ5utsKWWj1ZxTSWEBSk8+isaKco9qomkR23xFesoW659dvDlurj64dMJld5JO
+hZ+CWi0kQxeIcLQ29jpHmW25NjVDvXtmi4RJSKQxAYAUAkcvHJG9+At3RpT+Q3CKI6kbAS7BO+e
SU56fzYvLbbaVh+gBakKlpxyxSTd10+G320+yIXE4aP3gmyeLhdE8ygs3pV99QEOUd8aeYZ2VrYt
RA8s5Ho6SQyWTtWoDp7wvFMV8mFaV64fYYRGcMco4ujRYczDL/ZMWdLuKze1Vfb7x0sdDVMZ4n3T
OY8AKbQonw9jGdllrRIRVhsC+HTn0vK6tFF7MScxjiNWuhyfsWcwWCTlVtkt2QvK5ikPbaU3taap
Kb3+CY7eMwUGI3+8tHyiRIE/fW5zJ+2GphZIQfTFZ7Evg7GiXnHqXRuxpHXJVCngSOm9ZcLeZAye
vCJ4qGvrt/7MCQyXoLBbfr0a3tOglcregHGOPDImR016Q9xf6w9quJsjfnADMvMTgtQDIEo7IYBw
pAn7MXXUbX6FNThFkqdxejcr+wzxFqvXIReQtpv88W5l+3jj2vQaM1bt+jcZfvVIHf/MCX2ILWY8
rKqJlusnK4YbaaTELMplTG1BUU+SCtTNlWUKik1JXZfHspRmaDhsqUdHZ7wdMs2f9gcnH84PkhLx
RzHxqe02ZsWID6JYzZ72GCgLMho4CCkFjg0pWyIsgGdN3Zpeh3yUAY6V981Ha00UgoAu/zUOovcs
a9ZcItlEAHYopDLDEG7I75bDCMcbfXA6+Js9LRPsdnbNcu0Vohlivv7saxnciHBsAt1CK/3MlW5O
In2ras8t4uB+i2KlNYEP1CAke9aHphHajxEOJC9aet65qXc4hjq7ww3UOCn5lhOFbrNXG+v25AkG
SF2jae4SkO9E8zvGu/Y31ZnZpB8vVkOHGGtRu5hg/xfjDCtdAKqdOH9cnGvbeJ1e8HcrPsuaFLvL
UaRLCQIVK2O334yImV+U1GGObJARAJ9ZsgEzvC5srcetZuorPMR40iOXDtcsCZX6Se9mstzA6Beu
wY55rx5kyJ7vvPNOqf7SmRVAsjBK6DI9pbKen/duByJyCxAtqukl8KguBqQ7U1f8HMbacsOrMUZe
yfqMjwr8yTTamB6HiAjbTscVnvKVDHixOEm65RfZB4NPXEOEKv4M4yjzDYWq9UZExAirWtH7TNIm
SObAgLe0O27wh5x06fZ/n6n6FyYtV3uu45VqN8nNYrA7bHXGcfD/CR298pzfa0bXsacIBj8uiBii
9VDHJjLF2aUTgOG9ZApYrEu90dNDsX+Om8eG9oJ67MLNpkyJPvQV0/6EZce04uyPTpPuQ3ZYCYqf
J8KMmcf6n+p/Ng0GyOaIY5Z+qwrD/e8kLE9jazTBd0AoHeRbsgY6LFuD8N5nz3jW/AfkCgIxbzBs
xzLDCHE4++Y7PFmYx+5FcH5mpQEqRdURHP9qP8q7n6emKrCpRE1ruQ/HnVIW4PQIL6nHPjha1XQ+
Dt2U2Cdj8ml+3xERKskI5uXe3nG4siBKGAqJOR6f5XiW6Y8ct4f3CUxGnf4/KFy7cmvJwc2g1CMk
2b9PhpH1T8eKGRRif9ccmhaGmZLyRXV5pze61KXVYHmEpyDhmBH9GOUkefWeCzTSJH5Mq5aQ5eru
WJpybWNzEsg42OWr7/a6Kq87DwtM1hCDWCzvaE6CegsreD3wiCidj63wwYqwGj7qijcvzoKeiHiz
0y676z3mXIVwrq8glxHACR7zrjIMKgrRR+dC2hzpaETlNnbzE+wYRtanqWkS05I+SC+xmsTSNfvy
MWkJJ758ZjjKDL4KwDIrlnsEloDUvvN6nxHKBDA18GM6j9Zw2esIpMyN6QlRSOjWMBQkH0MgN+Fx
x6AGOtXJclRUcI7KfiVSA3xwsM4zLQ8yL4uMDquB16KKizucf1TzvQ1gSQXpvwD4TcT0/ncGbsJc
j4Tobm6n1jQXP03bqIriK1ZbTTXBDL+TCd32zloMMmYRsd8AK1k7F0DCvDSaR0s9BRQlYcE2f5Ls
f2Ayduzbuw/vi7BBVWB9N83rpNrrm7xwEJ/LoikpyL/+FwBHkAy8KXslg+4/3tFIrt4+OLjrRP7x
qMbdVM4s81k+ARXSGNc5xOo6DfcEQhZ4vJbcTpEQGJy1AAF+9B/cAoUjPb+OwDpdx/NxfwZcwvCx
1mAPj9J9uoiS7m/fbbhmOZgGT0rwDL0xVK4qsePUQa2laXQYObXuElKobACvkMxZPLHDxNtjhr5M
ryriGN3mfACYTyqRJlkJCbN/3CXI5dPapo6MjOXTWOyxcsVAHGM8QaQ6VvDmhWcTGeX67BGmje8w
Uq8LxBCjqRxFxQtqWbHePeqA6LaJ/u57EMO1Jkcpyopv8dFXZgnfMpDYTLzptxfS2L9FKj8p0Hqz
Zjg45JVd2oYICu995NkcBv1UjYdCjG/cFTok+JVCUdr7HLWa+zikNrlkFAeboCU0NiKxY0lgD2Kj
KGmOZIkarjVTMwYMvBPo6rYoCDgSRB9wDRZ66zp18RyDeewsNm6Faodb14frwC4iU1LzC2AXsyoY
ddfu6KvVIuIfsxxizbAZpGl0rcG1brQSGA32L/CB23kSAl2unAlZha5B/xjWsEgz0H1EBLLkExtY
h0T5pyqH4iTHXhbf57uoCLfS6OTzEi4NR6W4TmTa1POjivpFbXKYUgAMfQHxOfOyzjK554SVXOIi
6+3WfKvHiSvsh5e67cq/LCue4NnqlHqcfAGEPtNHPjJ67Sx4QtMVrWefzEhYOfY5hsvkfUpQzzWi
zAoF5vh8f9OWyd+ew930nCVgfaVe/9bK79cxhJuhb6U/PwxjpgVnf2GKxDhfgu+wGJqvaGIkt2c0
Xf/7XOOMLD3EdasmUEHxZlvTC7eiBuZRLkZ55xXpR5bfnDX1FbCn/H07B8EUlW2kOUue49b08l9V
Z9p8us4zA4Bfs8nGskSz0NtZAD4NlwZlbysa4Gm0BxyXIacX5UZaDQYC/HrXwYBoZbHigYe052bg
VhAKELLKtL26n6E5Eq4MTtS7hhgyrMnuXbtGDM7+xrbxmoaWYfI+FCrbiErCLK9LZ+eA4kN/fuAh
tTRJdJPZNThhX/D2+VFH2UhZJRBpAMsYBgif/yZM5+z1t/VUI7iR9aFtFV4S0KHTV6RS7gbrM2GS
PvpwPm4d5vaOGm5O3pVlKZqQr+856Ol8voOLkiNpE1SBRWnABrlhu0QBwIDjPQkUjn+13sxR/OHs
3vrtgLKsdxqA9ftlnhPo/q3EOw3PnJG35NraPk8G6mxsnB7mmGPiRPgcYA7uSEaULA4gIRfk05iC
KFjZWJH4XmeKOa1+NSiMwkTyADw2GjvzRVLqyBTW9CyovuPoRLten96EhjKne1rVLPSMRy0rkGqs
hli5Nd6ph8JyD3SHNGcM3eNt7mLi8a37HfSZQ6TAAmSfaZidGv77+8arPe2HG1BS2q3RyQviOAa/
r5SYf9I+XsYKH7YQbAdOqpuytkTAzqODtYOnxSmRgk+l47ycQBc5OEA28geV8WBf3mGn+70GlC5w
3fOYITrSLgWsfr1OAISASrlLAZxYkkWqlhOpIQBBgql5PTSed3W1DW2ewRPgNMirdtRWzIvO7O+w
vOyxwujq12ljkO01Q2iUUKfNAlhcRpdFt3a1VOUOveQ6K6MJhZOwtucoiuzuo/ANoTRYnUlByjJq
hPORbAUYGadCcgIGhyaJR2JzKm+9XihkujriOBYyDJ5PGY0U+KBN/ZbcFLFYUxZQN54UxHanCmH2
AKDoExf5N8lroAp/2IzitSE46rYSZx2nC1MS3nC9lYYal1P65nS4onIyqcqFeQ5eEp5sBOcO5K1M
3MC0s0N7TuBXAfSThGTnrBMlYtbfYuKq7uo8k0i5OeZGu6PQQsEOv8B6zDUljO1Fuj1aYZX0ORvn
48ZzYM6WTWErO4rrv7uomO4Kd0eZjkclv7Ie6j28hWapz4VhLOaryTboG0J7mXsSGJfJANbuZXiz
XBUGc6ztTDTeD70FxXlfpriYdLR1iXmoSt/k7DcvmnBBR4lwgwKUpKT+SdEms7ZxMJP+6pvUtsek
ORutLlangK5n31DQqDRQib4EpEXY1b6TRJQcVGO2f6Z6A+Y670cciC+DgPz5C8+cd/9PKCzjANdY
EPYgY8elxGcNdyZWbD2eNwMCqfKZEIos4gtcchKY9w5LuDyhfTvA//7l+b1JgekzKMwD8YdwNCU0
zWWErQwj32HbfvrQbqknqfNs0bZ3g3uVGcYOW2EkMqdSFauv8lFU9PBsdfic4z2QazTV+1btgdyT
WRkI+L+gpy8xecULIxX/8Pz4b+YzdZWeIHEHMNnu0DIllFthOsRd8SlzZGXvTOqJB+WhdbnWebqH
sopJeaPiq5QLRILmNs0ukGZWHq8wwlPZjxri/fwSKSMRuZZiZyFY1O0YrX+6wq8mvt9o4uH4VblP
3/8JONyXyfwExC+Bk9kuN7X+hMvCGHwPPaLawrm1Nug14EWJwO4mOvF4DOOVwiP/uwySu3VrWPe6
HFvyVhbtQpDFKWkWhpZMzBiJ+bIbPJV5inOWMmqHv2vuiaT56dEi9VtpFy2GV8g0MPN5K/Y5rHer
L+zc6G/Dd+A2TtdrJIHdP7eHk7FwuwdspZ7U7PHUmJasq4hSdjFW8RSPcfrJp0waQpyMbYrebbTY
DV1eHX4pqzlnuuzSMlZEajDE8LQ8KyIbShTKLB0jZ4gTgqqVWP4BcoOyDQbcbWCB58tYR63IFm74
1Z/iqeI6CXJLH24KrmaKNtr/6uo49qgMzflEaEuVN+9dej0LNJ8Xu8jpJrB8E6syqkQsMOn4EJqw
cmUuIFDf/SQqJH/3g0DeXvBr2zlAxQaaVLgp/5EhFdi/Bi8OyptlVTa5mZDkpT2/go/qPOhXfWht
fBi1IDyyasA43hLhGxhaPivIKx0kaYoU5+pOh60+tdPqpQLbrNd4bbQOJhKWO/QTEZkhZ1wA4CMR
HYcFvXj68IcPSVJCs/vao1xWHAjZ6HhFKgvbqyzWU9JJIUQWvZo/ECGRIYT50nnvoCAG52aA6kii
2Tnh4OiXqL5QgkMksqduBMLEBo33ktZzaLK4m98M6ZlsWvqhPd1nsR64eXSZo9ygzUn2Aic6Pwxe
krn0aTp+GsSAR8hyWMzHwh8Errh4pKZticPuyJOzEh+V5Fo2GfKM7V4iaFH1vaj/HE0LNIIpm4u2
M1HmEC0a1+IoKT1pCdtubjLWhF1CynarryvL9JjklYoqDU4jgkGzcth2j/M0i2VkmVjNAoSS7ChE
M79W4AdHb4WECXCa0KFXxD7nyS+WPfELzH9gGb1jkeNdLWRFtobDJqNLgettQbVwaHR0gO0vNlpi
8Ylgy1X2H87S3NXFbYzsqS89Mfeq2G7QL5dSDTcbchhSJYxR75+9er9IgSerDSxEzJgXkSRX3AUp
Vg/Ro/rgg+p9pQk+fXD8RqkjyVuKSe27N1O2+qpd9z58+wj/1brMMwsBKfGzPn5xUrPcFr2mwftK
lK9LVzUqhxPp2sXNDzL8g/gcQdnoBzNEisOnW03r93S5kSITGG2tyWg3HkDV2NX/lC3l+cGiGOqP
YKK0YizPUAjB3qfnItmh7uhFoWIfUHl4oNiEccvQUjbKgQpISPuL5IrgkOorj+DNht8wZvvi+fb2
8grK7s51NVpYCRA9sQC2Mm9S9t1nFcKnLy2/iNaBOllGiBRC5IMCRFRtyKQyJCkpndWW1XKrUq1K
lKXFOsNhD17pYvDb2MKfisRQS+3V7D2wpC84qlPlmsaC+NN2eO/B48tMp6FYLm/3SO9ncbyhqwNx
QFFfasKM5nHTOlBhssfQTvLpXcRckaF2UkctGm8cVe9h1u+G9aUMRXnbTVoqH6TjBpn8l69aQLt9
GkN7E5HKkR2BmoPEHr+Bt0HfD3L5+JIPhxpn4oTyyFXaG5Usq9oB+dz5FzmSuAhgjTvJ6x10UvCj
itE3dKI6RurZZLnUTPQPZIh1Q0dqLcYa2+QE75tpGPfNrzP91eRpDBIYLT73Sk0bNL1xU/ucnkHd
2Wdb4MKWIljLBWf1Haw5ugfaQLCWW/O73RzJNqvefRsarZMTGfyhL/Ow7lCa1zoFcboUwY6JtMZ5
gvq7/r00l2FoiHZc5xHitM5mwybVS865GVioyGFt6k1ek+w9qxo0AvdAvBb7U6i/OkyIEYX0rw0C
eww6qo0Fef0OOCOogq+WqCVWOane6ReoVxeydLkATKJtIaXb52m7C3ZM4ZFZQv5XumQ/URBkhD+L
754l3XF3o8hA5ONR7JYSTiqctNX+7LA7B6ue/wfRibwlUc32A006sb3uqvMwmGMm/qG+V9lDddlN
Cd5DMW8yV55LLp12r3Bh9CKeQEbfMKIqhxPyXyWiiy+AOBqS/KMZoUxMONq9wjtpyHXiSzucnlkW
a9TasNTQFzrqFrE6mWFNpHeBsOCaAQBpS9MS0GfGpAV0YUQXjrU0ynpDOZBryBdulmx0kuFOHPnD
Ijfxtxp6c2Vjds++TtV8iKdkxQGbh+hVQtpGfaH2HN0hNq5ozW5LVg5IFOTOTr6o7ghrAqv47Q0S
vSPTK/Zlv1sktE+vt2Z2UOMpwFULDiZv6k8oZeSHbtuE6yC6S2OrDJoDWzEndaDOiEthXxAnpj/D
FnFzPxQ7whn76agSMbgiLzHDZ7sGWL9LEtENIKe6zcgo8X+OZOJgIpGvzI738+Wcn882tq22rO5g
pqnoR/onoINW6vyXF6ACuvevGaqCSqIKz67dfkxFtenB2GJenSz7O7RaPQduCkjAjg126M/2tOT0
ZdIDp4hoEfWrPY5QTt2q0co3YUjkBhjQTXWyR3K3c7CRUj4qxktLaPvK5ntxUFPgXmvGAiuc6AQ0
KenlnLZrNKzzgJsu4Y5C6Y3YvA95Nc4sgazvSE99aEUPgl8V6CXruC5qJZrFaTKrqgzczVuV1rS3
3y7GNW66K4jdFNea9AFVR5FF8WQOHTlQ4rx9IDSvM50qC4QmOS30uQKTiSW98rCFXS87VsCySAPt
ymFS1RCMxfAKlz14926rrtKNTuHPBaiZFdX1eszRpvjTofZBpjudESTcO0qRAfxNse/E9h0JFNmA
BaQYqc+3ofLFy0v0YZlud89/hn6qO5acj8YXGWwtgceBIqSXOd2oqFCBRFg+Sww0Ze09j6X61lvu
oqKHWKSAdepb5CRgb8okQU8s9uN8CJ4TBSUsBoCYR9m3eIqMr2BEojeQHMd4gSCqMDTqPzqo1MpK
QDyx2WoF8PXE0gjusNgRW7Bq1Q3n+W+f2GK+VNiCbIPdJXE+cG0KiGmLPI2ssTKec2vuCR0JZPUb
XN2jiGAXo65+IeXxhDKKa/qhjNJ8jcTNztwZpOLmQ1tVPJAhBwOHBdsqRxS0p22K7bCj1JXLWUJ0
nX6GEWvHqJyuXb/XokP0SnNgvXVH/H8kcMB/BF+8pb7j8M+eGR3FfjQa/dYS4XQXecPNzRlLD95O
F6LetJ2/qgckN2duzweG5DdiiTlupje5oF/jOpbHxiepcJRT6riv8xTZDyB/X8mtWbEEnizsg76w
DY4k5g1h8O9rFvaeq0afyo7WizBDt0rTC2kl4/8bh0VW9sPIcOCw2aFzr9Cz/FSudPUV8fXeDyWe
GpjAC7SDdAubo8ia1qXAKhfY1H/7ZR8MNC00+nUogIFLYbvqN11JJJLsfDyUBwJ9dMrsBuPNtKqp
EtIj8i3MslMv504tS4yy2ZSHhMPVbMkCMJWa6wMJS4VezBB0m5BhEt9YoaQNeG+fm1Q8p03TFySI
YiTAV3SEyXFVlUN2/KnAzhfMc7YAE2Up7yVZxUvca1nc4P3DCYx0Z+ZICf5dM/Ah0gRbGnOsbQD1
iPBR5oFtklSXHPVA32YjKRPYtKxBAVieO4R8AXGbXznghE1EQg5GcJSY9GtU7DwR9t+/HklGcyMj
cpLN02QNit/QnumC0U/TB2qDSYXB0cblngStKG0orN251bByaoFitktFvYTIRcpUvb3g7TlzzLrQ
u+OvRF0aMVRe68qwaLTva3oT4oM04x1101nR9OE2x/REcRwYUN1Gi+fi157RgIff8Xr2UT3xSXn1
1q5fewCRwJX97CUytMdD/vfwVhEocVGH+4VbU/1RA5YWlLSvmDC+3EkQ2ZESiynCCtBkXf7iTudQ
9OrDPzF9vYBtcp83tj/CfcaO6tSIT3LDKEFecdlGqpJhfDLPd9nVzlHj8R5RYvTqS50RKmuJvw3z
z4cc3FRlZgKu3Bjpd/7qLvrqp7YLRchTNnCSoIoyq+7NQRCLxxG7obm0oK2hcg7Id/IxY9PlnwWY
3o9zjg0LAxREPW2wUYeNMyUREydfzeCCY59F3Ro9xgUiCvZY97zPRnou3SCwJj95+4h9ezry23R7
TZ6brDKNrFnZAqKw27V9pW4rtQrVfERSjLXiBNOYDC9+0C+SKSF2NkhYBRYjs2PEnDeusTtGivOH
7YfF+tsPtKV0jzlgzG9vjVplTyvhuCkzW9AKiYHQ35rRl3TJvpfeXKJfHAsX6ld72z8AAvD9BXNb
WZaovLzl12q/XbQtDGKgHPDa0c7zfH6iBxeFQLVd4t/+ka5ZQRR1jCfVG5Gcdy/m8jTR330uloL8
AHgnmD1q5cOGHTKvOaG6rnf11apjmh3K4gAlm08Yavi5c7MTOkCplw4izfJ+8LKyHWu5G12uHmSJ
fn/PeWq6yEimStJQkAAhWUsLXIdYwmsP8mwFDf2ruQEsxr82CqzoWjL3YWf5QG2B+2xwwSdn5ghG
v/LNOyCqFEiS4Jw4IjfQIglThU28S2pKQnxiP/QJBNkM3iR3dgGcUIf6mZstqIq2yYxlWTqTTbxL
px0ZdR16XWaWI1mBxdz175Ow27jpUChwPsEgDtDyCDVE1MNk4kU9wG1FZW/ZorzLDx+6lHEt1u0C
Ujzlc4NaRTfVPW9mF08EckmhNmO6l9BiW7ejB4hU3DzSAnbFG0PF+JOq1wiG3LPCf+P2XXhL/exq
sBJtgOv9Fc6AnreYCQa7crkejP1xkBBWk9Js7Eas4BQG/Fki/QfNf0+yd+TyTvlX4h8EvYhR73PH
ZQq5jqT1WiFab1hg3hb1CQ1zExMvXJp1DIhKm8W9nhxZ50ziF0sMsI0PhCiIqa+0rYf8gpOTt0x2
XcWwaCLINsJPFZlSQ1c04gXYxa7jGNQ8wfzEVhWoFqniZcDUhrbYKUDijCp7hQXamcR5jdW4Feud
LV1YDn/d9VW9h4QvYdEueYSVtElLi99Q9/TDFxXiQ1zbXFP++NDqTwoqJLqfxZ33ows2ugs/rl4E
8O+BWEhca/jHinXzhbILM3OGmsWUP7awnioolHhBWJH2UrE8sSdHe5vDUyvVwr1t9UXWlMN2WmDq
zolNWXiIIiKsAlIZa9FEMeKbCQ7l3yzYvxLCpUagefKJB5XJyA8EnbF6xv6pJruP7QVD+aIz4RiF
wIy7FImHHOjBkjpO5/DJY6XiCbKKZrmEPUM7CJPm+mbdjnZcAn9V2s2kOjN76HY/ADaIYCYkmTIb
qDf5k3biT0hU+NLYZK9vJKuhBwEGUvL9STAfTrjkyVuhjQYV76rbbvPLoak5fYvVO9Y2Z4Is6lxm
nxo/B1WL9K73rGBbihqPwGYEV1XLu9YxvRvwSkbITrjGWDbNDVwXEMOY19R3ZfDINHzPhXV5HGni
LYfYM1ViFIFcB2OT+bfT/WaAdNkbvWI/ktlqvxBODxk3Kn1SUKiEojnehB88BGwxz6FJbkZfH80D
GfLLBJu3eXozpBTiVh1rQmEMJkUy4japnJCZM70I3yD+PjCQLdWBE315+6J/94eQytrF0LXg1Tgs
QAcQby8y0jJurj8IEQpf8E7GMusC/el4DUl17ebmjicyAQ/11XzVO05k8QZ8Xj0D+KhbMw558pAy
8BjJ1nURAcXAGC5Ci+rPfZSavM6WWZb/GUVfV2gy/qzrnQu4S7P+FZSjvTsIk9QN2uIHtvm1NEyE
mktt03rnpGVOCxYGksVYCIGSJTw6ZzcPc6PKVaz3DEXxoQjplq3IfEDy78oVBpmzaAjHvjv4p+Fi
RJefV4R0sqmACi+Ja33ef66/t3CKJMBmxIdUkPtF3ZknNLBRUU5EeZxEdlLb95jGfGSKR/0gezbp
JI6Fx9zLt43RlyVhNHVDJrpi0t06g+7MbXpsLVcJCtJ8OosvP1SYsHub+c+ltHgSSXSVUPfcY550
Q9Q+bnG1CO6jIQeIjYKVxw+/xnhUExHniAl5HZXZ2Zp/3rWvaajztL3o6GBbOIsK1484GvrxuVTZ
uQ7oTYxzyYwdMkxWLuPefw3xTAumkCAembGMN0VnoCBdWLjS01fW6aEQ2S1dmt+c6FlXiHW0L8gS
E0/CSReZr7RRzuwYiChuSkcdYshwFF/ORabjC6vzsHfoD5pgujuLLgw+kbZBOkL9Y1zJVlcehguS
niVuoKMibaL7J+1dYOHBtoerfBvBpd/3CbyQ80+wXzxFlvl6dpKZDNxubpgmG1sdFBOH1UEhjMln
K2yNQeqQ3uJbc+fOiAskFHni0oCpNGJwC4epN8nQGaR7cH5IbE5+jamauxW1oodOQnb7X/6CNUZU
T3YaNCM8IX+SOMlcasMgkeZBP9fCpSY5nGuFkjez1i9THJEAD8HXTZ1T958eii8OqQbnVYYFm1Z8
T+L/NrmMCGgnqNdcHKpRdB0JliEs++O1x5PSDZUYjf36vxLZs2UGGajipjuXLIdhztuIxhVIhY4F
Oak3Unox+14LJJLL21MLwD4dT33OZU90oNeMSI9kT+t29PKisA4ZZ2rojU3BdPuwmMLvYNevsHbT
mqKIAZ3/ExhJqJ/o5ybQhK3DHQrPZ2ZOjgdPRIPEArcWF9irkKWhdAS0VQkrYkKptE66UaXQjwAX
tsOC8O96C8J+DkIl9BVDdtkIVps6jKWuZHwCLr21pB2WYy3SxYalByQ7KgGkSm6+s97oDOd47S0l
ZmCoUCo66wazWKvRfDRb3sSfg898jevcFQNafhkRr2lXdV/pygj6uGVzfowMckv8wq6mMHU8ou4A
6FCT2MYB35jEgdU7x/lofhTktREnZN/pfSSTJiU0OzZ+v4ymcQFfuzzUC+vNDAE4n1BycrreRQ0y
fkmfHacwsLOdfxjrOxQiwPybt85I1If/g/JI8a2xxa5pT51qrMFDPrjqiPzHncuYylyhlCn5PNoj
b1stCa9MdMADTjq6Jt4dee+s2Kh1awyTfn7jBzalMcQ/YPiGRBZ9Hj/BVWzv9ixQ4GDB3jVGn9R7
r0JuYZQGk04eGJsdRnEsbgrgoSnW7jUHBTuS71A4VDCQJyn8f3ZdTQO1tc5ljoD8xOxPWSbpy3Iu
cB5QCqbQLFa2TNEpQYF6lGv2nvWMzX7dSpOR6IC5pRUqq9TIJd6/87HTUUojPjuF88YOiLLbEz9v
3wVxFB9Wp2NeAxwsyOboFnzvvgDgjKIPIigVLqC83DjeN5Sf+sGSCx/ZcNNHiWuOfwg+FxUqak/A
mhXt70IB84El74U5FP1yPEVPFBydCi6EECsSy7JDZ7sI1Md9cftU4euFRpzt7YppU8K5VraDMmsS
H5EOE1rLXoFOxa4Zr/XoGmX7Vxs21uknrmjuSf4J1AejE5xJVkiyXpclNk2kH7nNMMy5pvaJ6dfc
On2iqHZ4VZ9ttU68Z7jA6quTRCRqTwklEMvqIYccbWy9pbqoe7xWHDYuco2Q3Ei8VqYpuvbwPge8
c0VvrWnlGQz27Au+k8jO2616pZRjxlfR0IAWpkQB3b9LhaxRYxNKgkPeArmDs04gDSIkB7oXFRkx
KeSlHQCVXcUczHDg52+6bLSddWupl3HL21VqU4zEXaq9IFwYWJv7iop5EyjuMN3dUL/uC1zgIc81
fffU7E5TS9cl7mVOEjQZDCyTT/TfV1y7fh/Sl+Y0VJJ1iMSxdMNm6nfjR0sySCnKbrkSmY7PHYke
KuEUvf+heV8Lb+2ieg4xr4GABj+vK2LPvLpxSJMRH/vHg1Py08hKbbZg/VK+Ch/HYq7IJWzqqhnS
d2faEUmcloowFF2CiO6yM02R1tgsWoUiFSvzhAT/Do/FUQ3+qoA17Uzmb5dZIAP19T+551q87BML
5hoZEKOpo2aosX++W/P+bSgvWczEYKLqwOf07CeR93ek8hkIEBLPfmudN6+zRMEEAY1jE34uIcOi
c/r+3wJc6uT/R1YobQ0IihCNSvPd8EsE/a2taTrwU5uxqojlM51S/79A1RU2jtBgyDOLGcA14zso
ZduPwhlTdTFCVB4YVR5B4fwBTb6wVB76C9DRtMlM6zaZCbVdBEGioduv4ZegZYshuq79v4ncC49j
Bace/x7oNN/pkllixuOMiq82ACisjoay8qZFXDcfakbJG61VlrOSIl/1iLpteG6Rrq26P/y9ookS
Li0kwP6RjordlVmtyGeTA7QzovheNEW7FWkEP+mzCsarKmdIBIA3EFPssShsL4kOC2Ozoo01PSoe
Y1+GPOWf+R7gyZ6TXC6vBW0CmHNFy+SAx8XQz7AXG7XOInkhdzAeRpeQGxhL4yh4ld1Rv48HICKT
5puDtCrn2tkuPAHGhk7xpQTK4DmJYLY+nlaxlrRvs2+qKzh3+lq8EHXktwVkTvjOYUQZBotK7TpH
hBBNEn9vJi5+f8X8/Et0C/1gVJ0SaWb+L2Y0yWx9KExS2tOCMARZn3EPtrhVz1dANprw67BTtakA
Kkbg26f7bpRFb0ueiHtcR3l00qf+A8EYuR4NVEI89TF+X5FVJzoQbL072Lme4feAt+ex4S0niAtQ
mQyVi/u4ZG99PcvPXi6cFhlr8mCvk6e8VqlsclAAO1J7iQ6RbIhM+TTIrWaK9B8pSyvwSkOdxTzq
R7t/8+lAFg+Ct7n+Om0gbs5U2VyE18ArnfNCgjCqoZCT4se/vvP2HZ5iXls1+CKCgRdXJvi5z/oN
vguDHCY/kKJBnow/P56uXEBXJ3bAUromrwhO/4lkdX8OHK4q3q7CD6koKpGnrtOBmSYMJuBnILpe
+6cthLpGcR+R7sCgy4E3I53zUIfBl6vNz/40Bk5vJgXv24OVNMEo6ESkbAr4hROyIDUA/vg8XzIQ
ZFsghLpbUlT95jziup+WaMdOaiiB/NRgmgWiaioJCC7wPgGVx2KpI4I7XYca4L3gJ1eaYFkHFvXr
RsMnRuCVgQ5c1Gv5KKnwzQrevBos0ToanCqopLz4pAKiiBM14FR4uCa7X99+tcWvu/3moS3GsCxQ
VhxcdIWMGvS7yLGTYTSLDvSglyzBN2C7EYDxiYEgP7iAvXqZrEeH/24N90wmoz82xQzZgXdYXQ7m
cPTqDhQyk2WNj/lBbX0SYWdBeVGGHrGs9IVFMx/diGCyBhBkKJRVDf0lVJiECkGROM1SnaL4uqdK
jx10HKuxOsB4jJIDgbIm9DEPNY2i0FjRS5Pp8/XR7r/u9F/1WsrnwtuH7ZjWBzQZoRfpSRxV/HBp
XZPNaQ59m8B3KGFsdYLkFR9MyzheT2qCZFfOPZgOCOIWUbGN9Sqsj/igE6BAn05NfGve/yNxmqGZ
racdb/8NHJkvN4AKcglrkkOtMiE7rBjytDmgJagi/MXvvzPkaY3bTM+osKxtBTl8FOdN24mk38vJ
dl2dfS5dNTucx8kvpnn3vQMKBI9CXVPeY9AGph9HAtDINANOFa3vXt/mHKmkTYfYXty6Q1UeQAD9
z7m5xwU9zGcZvS7+BODMY0FfF95QS3giX3FfcBVh/964GtXKvet0BX9qCdLB9OIxGYoWRFNiTy/Y
mai088+9Tyt0cn4ujPMMl59pdSKnWwNLNcXQQvmbKajllr/jjb0kVyvhnQa6jLLW5xC/kdrOcZZY
R/eSqE7b95Mj8xWptxOVLY7tfIOhDlR58rRFc8W2ZGkhEjeTEPSMgqhdsrT9s9tT2wD+UAekReRy
YFUPGx9kNhJHlwNiZKCnDTP5SR80eyGkcnczs/8qBF9v+Sh8jvH+7hGv7jEdyvPKGTfYNdTq2fk3
Ihzny4OzZ+JoqKStAbWmNLRyuQlnOaf3IrfJhj+yu8U3Zk3s0R5FJlBSZbYIqBySEzye/6m0mXkj
pWvtQFLwpzdRrX9fDr2ZpI3d9AfZNlMlNhJxf09XuF8vKPNUBZmSRYYOQn3drm35X+lJsZUjuMXP
8R5N6QF7ClWYcoHUMkjy4L+6I8rjMlG9oL6NcODAeaHR3sUPmL1k1RjiYYhxKhMWKsXV8hU1BBOs
ne3WsiYUI5F+5LdCG2Px9NAR/NVxvcrmxOV13nsljbYWBgr/MWqQQytm3Pm9l7iDtpK4lO/BwtXg
8V0LeVsYD2PBEYrB//s/xzWtFJSmXzlqvNMubYrsdA8BQhXl74pCTXHK+QRbzyHT6hwnp/LI78C7
P57GTPZtKgfzdk/kAi/igQ7xwnEzT0J1uN/9FSGGwx/0UKx7F8PgiUwNKYcx0HgV+VRHkKKEb7Vj
KY4OMoVICIgefKbuAE/9Ny2MnmSI0P1a7Q29eWQdcOheNgx2g/jBkiNKpgUOSBWtTOoGM2hEvt2I
I3r97bBmrYquPVN4cEG5oXyFyvfQEvinAbRLaKTB8IWhVTHfDVbPklXq9gEJHw1Je/fUzRbFrMFB
67chfmK9ZGwUnCXhPNTDQs1CWtlAO5YPcajUbR+Dd6MIlU9KNxPjmyv8GW7lALu+f+VI3p6ZK8vk
+xZ9VBiTUja3EIxR6GyK0maJjhXqWJ8W639EA5/LhQPGWoSHrMcTyD6dHeAk5LqBcvPue3acltYi
NEM0NGLh404JSnM0wVj4CtAiQ0UUTN6/yOzrz/+DcrINE04llombf+j1PsFb5o0RTZ32LlWfQJgB
AeNWMTaRLYzn/tAFpU8zjX1HcfH3LEAxKD6goQ09IGh0B+ZExwyf/Yvn3TGjy+HOIFZoElyU8XMA
pzuUA8Ly9cvf73AghRnrkdiQJcNvmSWmFhRUaR2u3PYq4gciFMFjfWkUN5h5y7Tyar8lO9oHOYdK
mLB5Xxi6ohF09C5uEYqqH0weP3yMZ2TMqB3h2XvoNlVSaI98HB7yG3P6RhMsfagjlo8jmNfPBp8f
8oioH/qZEj5M2hwpqsW7u40pwZ5RnhMUTsIoy6o9vmY6dzC75XxijeEWh8UwQZyU3fWqljb3/D9a
v/LCHD3Gxk+feSfrxThL3O+52cWCDbgPHA6Nv4fw5rVT4YycHUd5tZixt31rwwSuMu0JmI20ROvs
1tR+AH4DrVBzt8zVw5Oait/L5pswk8aPk0P5V1sLyNOp5/lblJrhuRkbDvYfpziS3HV9P7fEtVTp
frix8V8uU5EIFtlq5ntH639KGJL8X8zzbCLSXm7Ir25wOfPmJ40AQdVqvT78rPj40YG65VJahQ2p
L+BWRGEgpI3ai/R8vnGQCVwqMoZ9dBnylPFukIy4J/FkfOsBH17LCPy0M8GA8dFHrMUCuWSQ2gF/
IKC3ZhQCKy7L4t+QkzcOqoMnDyDOs2ob1f6WJjYBloBwAVH7dt+yxW/ZqnwgspujKDRfhj8ttxCO
dZ6lWb8OqCi6y2FocB97wjg7T9A/fnwwskoYG6V2kelDzFRbiHDasqSEcVeiSSOaa8fwhpiRtkXN
7Et9PTxXWxDAK3Pw6tUrITX3+B4RCltWeYl9Ta8wYY9hS/5ETyPIrTjIFlrVVEYFKPYKABuDJjuA
U+A/8Pk9XINLdZOGUxr/D02f2J0G0bvjd0pbA1NEN7qmcHNjWxzGihqlSZpW+ZpshSB8945PPMgy
9epuA8+xJolbcGlaVZ+Rd/NmqAa3SwcYvXZ4sSXCnZV9Vmtv4yb8qsF6Eho4U+2mBQDcPmJhevaw
H2tubUEounsIZ8PPfk0DzOWyMJWeukVxR7MfVlUgdQD/8aBaXjxFEqlcbAS9q5Bdgx3oJpyygIWw
Tx02ydlVkO8Wnhi6DiXCBS4nOMwEoPdH5wwMFYaxiYkfTNeRjrfz9DZ5wHL1BHLHQLhE1YqhdpGu
KK/K+G94Wsn2j+q8jXMSTc4mLTzXrixqz0skenBjmd9tuINGWxn02qnCB4D12SMGqb5Z4nY2zSk6
XsGveeAcJBOevqVOHI+9mS7M9uOq1kh+GoyXZ/CcVSY+kpMMYUqOrR0EofjsrTTQUKyfdk7Y5psR
if64plPO7h+1ixFywpBoB2KNBngmxR/9R+FVSjN724HUl63hL1SnnNqcIlyd8Q5LbJ0SJmqMZVyS
O3w8BegiTGeC+Jvv4/jsqZqImKCceiPH0Yqo+xYiIXyHauCyZew2YIP85kntUamUIWSMLFu1U5A3
tkWWfMntbnsMVYkdBXGdvEHwfNt0uC90KeXIFlYT4JJLIeoyc+hSxc8nD+nsiLGA1rLlPTWb18/M
jQuEWMbfR3WHC5kPZ8qEVTIuRlCoRLee38X9+baQyGidyh/xNYFUUGOzWxVoXhKO33fXGXkhx0xR
rsHECJBTiO/8JrSgg2G+T2FD8sNzV7in+3ACAF6JEwYQTHdVX26K/d/FBRNAGUsD1HApfjnBsxww
sUvk6waidg0zTpVXO9hkGMOKRnZEfC9aUq/LkzQOZK7yAOvw61ETob/82+jeE1HweMdzj1mlTL6W
LaHrqqUU7rlwDLaiOzEeLwWJziCKu9/cW2FCFFPXOa3zFdmxTrPt0mipDkjVwjo/bl7bUotKBCA9
AI59i9PuSQSEcfMS+5WoF2wnFl2raPSXVHeWQ3zZKlIL8f+zVWDw6TAEzJ+TXSBd67SWFTzswS28
azsdvvmgA8WGkqqA8cAwkJShFp550mTVuD4584NbIVyvoCnFtTmcPU7OTLQMY6DdIkIFJ0Ple/cJ
kAnAdXxpa3UsFK6mttWO7VwmBFxaUcQHzbduilijom4gpvLTEIzDPeM6u6Ato1ALmtgh9So95Z9T
Pzo/JmkPnYfyjTLKw7AiCKn0/qWCTZVxcJXmnQsgO7yCmZ04u39hCtx6g2S9ygH2EReURvM5ijgo
crEcmJUCblaCI4vqjYBRexgRroUUGtPSXd8Jy8pR6ULJbMcGfl0S673qvN1TP2ztFwsMUipxKoHK
L8DM58NrUFDnJAYHc0Q8snbaWInSo/AawcwZjw3pJZC9nFhYYq1mDQprwUur/fg9aJfWUk7yByTe
hja9s6tVjXEP4YC/C1Rg6zzmxC9LZR1D+kqZRS3GqAUlFS/NvU/M1wIC9ezk5lNU2qu8Q1UOtZCm
RIPg+hj1tM38a7WyxV64tfBAvDkEh/lZ/0a6Oe0qBwg71mxhqqdaR97qrNoy7bQCr14mZXj/JcaJ
nkZwfv8alvPz3xGHv8VChaPf5JNQMt/5EdW5uxomQ408UJJXSD5VH0ziAljVwW59ZUYhKEM4/nRK
SLF/wWhg2y2yb09YUWFAdSeTcSmPCvxZ4fCGUL/gsoLm8SUFyp81lLKB2PVM1AxYY417b3jFVEcU
nBTFw0bIr7SYaba8TGmOLJEnpu6HGF18YvSpEGXYC+CtQWWEmiWZqAlWHajiX3PjVdUe+rAbtfTi
5/Q+2+M/4vMsN8BvZm7OJlzdHnu4CN3yTUgxV7ctl34crCRKsF1iUc+RHVh+jdLufAMJ6M0GyS6S
3yP4ARBN08Orb5RJWwbPajCJSCdzcDEyfbYzicQVF85LiQmCR06WizNAiHMUd8p4V9ZwO0Cm2K71
Ci8NQaPVBGSKFrh3xo0kXXhwM0mzyDTCJJltiTTgYgQ6+vyyo62LlECsYBwZSf2ccw3Vmb13xM7M
7nOmh3ATWg5dou0Fss7oTvzSJcX1xZJsUA4vHqF5AgahagG/9VVb2HXdNsDpMaL5C53Ug9lhsaGG
TlOC3MYi5mVzSkwm3urPEsF3FZNf9LarTKEgUpYqHsGTinKzDLbUTAfztV3KKiKmjw7S+UtD767l
4YVYfsoxvpFtIbQ+SsfUQC3ivy12uwvFTPmxb3cN2iA/soukl2baTndOd4cPnHayy8HFkNzzqO3l
Y3dxDk1J3AzgUI4BeCwsvtzv/8wm6NC67PTzwNJgSLoZzwo+7EhY5v39ze2CpV8wStrVhwNI39+h
BnqDk3rl/fHRMCNC72TODcYXn4k52Fe1csdH1U1u6M1c7WPKstEHbtpbVijdDnPniMbShX7mTwGC
be+PxlI7/dcevypP/ReAm99dkvqmvbTDpDVvSdHf8+LpJUM8UthGFAv5qcqrymhfncrq8u0GpXvK
FrkfCfKl6jO84avCzfeloNseeCH8MAHElpomRJIZsglJ+jx7lmc8v6wur7tLyJ6R8b+RQSgmyMog
oEDwXijBtaJpMhWO6B5FW+dCItZrBo0i7NisZU42TbD/ft/0j8nYeAx6KK4wePQNL9Hd5gayKJq6
w4L+zBxeey9D+0lGNZeSPZAB0h7wQiEdjkriXaAvKX4JqceRCCXsdkmjLDk6ZF9sFTXVKoGjoEOz
NxFQJ1nvLt/w95rFBQk8KxqojX+j4/xABwFXMsgj38YSR/zI+W7R7VYOVo1wJYixw2AIerGgZceY
rZK4xaoDX8iPJyF8x0txnEq6fenQqqDQOZcGEuI2PREEdC6wn+fLNqhyPTzuABwpLBWOQXe34cgq
rB8EP+UPx1AnqqrMQFZzhqMTBxRx+rQ+bBPCNO2Nw1pdv2tvse5VAeP3m6YDJ991iAHCRjbnPX5p
4zKYSGIEf4SHo3Dq4e4WPpWkhaHKvh/g5X08oGM7C3TcGkmJD2AbXPnF3a5V9Cl461ZQ+c3bp1uM
oQs+3mL/dEKMLyGu8Gi30Xz7/3sZiMlXkm8aMyg/js2NKK2BR9eycm1I5rWEJ5ij0dJA+DhGjkRy
BX5ucmTwqS8mzkajbpOL5MwcYX4vJg8TWCrkA+V66MgRvlueLcgX+SuzAfgcS63+CfVruo6AwO5v
qQzjmv6aZFSisxeGRVUccGsKcrB3+aWWB/2+MxMcxhZc+0ahaV0JwdVHqHfiJDB83I62y6Y4E46K
ISBcyt4MkX/7l3o+EWN2q5dXzJVm0TDogQcK88ggjbUHq7id6Xy6DEJy5bLaSYj72qT5k559JLak
5zjkgCdvQb/p04PpjPtGJWB3bMR+EP9zPk+uLwe7XsJ7mbKX6Hakb5S7kAxE3YOSmRdoaBZc3dd0
tvSq8ZAe2Y17jiL1GglTiIwROrZVpaywg1+ChSO54vaiqtySEYUR4518ljvj4edLXFe1Noh5NNrl
MGzCNPnOL0MKxi84FZddzE9K2eI0/KZcmmRhSssqmWb0mDaKbl2bV+UZCqPpAYS9ehnjG1pyaC24
k7bWFpYKWX/owHAA+8mr+m7oUpNCL1N8YZKJ3n5pg63ukbhASg==
`protect end_protected
